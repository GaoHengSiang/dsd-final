module decoder(

);


endmodule