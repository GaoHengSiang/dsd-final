module decompressor(
    input  [15:0] inst_compressed,
    output [31:0] inst
);
    
endmodule
