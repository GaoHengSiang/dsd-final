module mul_unit #(
    parameter WIDTH = 32
    )(
    input             clk,
    input             rst_n,
    input [WIDTH-1:0] a,
    input [WIDTH-1:0] b,
    output [WIDTH-1:0] c
);

    
    reg [2*WIDTH-1:0] z0_r, z1_r;
    wire [2*WIDTH-1:0] z0_w, z1_w;

    dadda u0(a, b, z0_w, z1_w);
    reg [2*WIDTH-1:0] c_64_r;
    wire [2*WIDTH-1:0] c_64_w;
    wire [2*WIDTH-1:0] dummy;

    assign c_64_w = z0_r;
    assign dummy = a * b;
    // assign c = c_64_r[WIDTH-1:0];
    assign c = c_64_r;
    always @(posedge clk) begin
        if (!rst_n) begin
            z0_r <= 0;
            z1_r <= 0;
            c_64_r <= 0;
        end else begin
            z0_r <= dummy;
            z1_r <= z1_w;
            c_64_r <= c_64_w;
        end
    end
endmodule
module dadda
(
  input  [31 : 0] x,
  input   [31 : 0] y,
  output  [63 : 0] z0,
  output  [63 : 0] z1
);

  wire [31 : 0] P [0 : 31];

  wire [929 : 0] S;
  wire [929 : 0] C;

  assign P[0][0] = x[0] & y[0];
  assign P[0][1] = x[0] & y[1];
  assign P[0][2] = x[0] & y[2];
  assign P[0][3] = x[0] & y[3];
  assign P[0][4] = x[0] & y[4];
  assign P[0][5] = x[0] & y[5];
  assign P[0][6] = x[0] & y[6];
  assign P[0][7] = x[0] & y[7];
  assign P[0][8] = x[0] & y[8];
  assign P[0][9] = x[0] & y[9];
  assign P[0][10] = x[0] & y[10];
  assign P[0][11] = x[0] & y[11];
  assign P[0][12] = x[0] & y[12];
  assign P[0][13] = x[0] & y[13];
  assign P[0][14] = x[0] & y[14];
  assign P[0][15] = x[0] & y[15];
  assign P[0][16] = x[0] & y[16];
  assign P[0][17] = x[0] & y[17];
  assign P[0][18] = x[0] & y[18];
  assign P[0][19] = x[0] & y[19];
  assign P[0][20] = x[0] & y[20];
  assign P[0][21] = x[0] & y[21];
  assign P[0][22] = x[0] & y[22];
  assign P[0][23] = x[0] & y[23];
  assign P[0][24] = x[0] & y[24];
  assign P[0][25] = x[0] & y[25];
  assign P[0][26] = x[0] & y[26];
  assign P[0][27] = x[0] & y[27];
  assign P[0][28] = x[0] & y[28];
  assign P[0][29] = x[0] & y[29];
  assign P[0][30] = x[0] & y[30];
  assign P[0][31] = x[0] & y[31];
  assign P[1][0] = x[1] & y[0];
  assign P[1][1] = x[1] & y[1];
  assign P[1][2] = x[1] & y[2];
  assign P[1][3] = x[1] & y[3];
  assign P[1][4] = x[1] & y[4];
  assign P[1][5] = x[1] & y[5];
  assign P[1][6] = x[1] & y[6];
  assign P[1][7] = x[1] & y[7];
  assign P[1][8] = x[1] & y[8];
  assign P[1][9] = x[1] & y[9];
  assign P[1][10] = x[1] & y[10];
  assign P[1][11] = x[1] & y[11];
  assign P[1][12] = x[1] & y[12];
  assign P[1][13] = x[1] & y[13];
  assign P[1][14] = x[1] & y[14];
  assign P[1][15] = x[1] & y[15];
  assign P[1][16] = x[1] & y[16];
  assign P[1][17] = x[1] & y[17];
  assign P[1][18] = x[1] & y[18];
  assign P[1][19] = x[1] & y[19];
  assign P[1][20] = x[1] & y[20];
  assign P[1][21] = x[1] & y[21];
  assign P[1][22] = x[1] & y[22];
  assign P[1][23] = x[1] & y[23];
  assign P[1][24] = x[1] & y[24];
  assign P[1][25] = x[1] & y[25];
  assign P[1][26] = x[1] & y[26];
  assign P[1][27] = x[1] & y[27];
  assign P[1][28] = x[1] & y[28];
  assign P[1][29] = x[1] & y[29];
  assign P[1][30] = x[1] & y[30];
  assign P[1][31] = x[1] & y[31];
  assign P[2][0] = x[2] & y[0];
  assign P[2][1] = x[2] & y[1];
  assign P[2][2] = x[2] & y[2];
  assign P[2][3] = x[2] & y[3];
  assign P[2][4] = x[2] & y[4];
  assign P[2][5] = x[2] & y[5];
  assign P[2][6] = x[2] & y[6];
  assign P[2][7] = x[2] & y[7];
  assign P[2][8] = x[2] & y[8];
  assign P[2][9] = x[2] & y[9];
  assign P[2][10] = x[2] & y[10];
  assign P[2][11] = x[2] & y[11];
  assign P[2][12] = x[2] & y[12];
  assign P[2][13] = x[2] & y[13];
  assign P[2][14] = x[2] & y[14];
  assign P[2][15] = x[2] & y[15];
  assign P[2][16] = x[2] & y[16];
  assign P[2][17] = x[2] & y[17];
  assign P[2][18] = x[2] & y[18];
  assign P[2][19] = x[2] & y[19];
  assign P[2][20] = x[2] & y[20];
  assign P[2][21] = x[2] & y[21];
  assign P[2][22] = x[2] & y[22];
  assign P[2][23] = x[2] & y[23];
  assign P[2][24] = x[2] & y[24];
  assign P[2][25] = x[2] & y[25];
  assign P[2][26] = x[2] & y[26];
  assign P[2][27] = x[2] & y[27];
  assign P[2][28] = x[2] & y[28];
  assign P[2][29] = x[2] & y[29];
  assign P[2][30] = x[2] & y[30];
  assign P[2][31] = x[2] & y[31];
  assign P[3][0] = x[3] & y[0];
  assign P[3][1] = x[3] & y[1];
  assign P[3][2] = x[3] & y[2];
  assign P[3][3] = x[3] & y[3];
  assign P[3][4] = x[3] & y[4];
  assign P[3][5] = x[3] & y[5];
  assign P[3][6] = x[3] & y[6];
  assign P[3][7] = x[3] & y[7];
  assign P[3][8] = x[3] & y[8];
  assign P[3][9] = x[3] & y[9];
  assign P[3][10] = x[3] & y[10];
  assign P[3][11] = x[3] & y[11];
  assign P[3][12] = x[3] & y[12];
  assign P[3][13] = x[3] & y[13];
  assign P[3][14] = x[3] & y[14];
  assign P[3][15] = x[3] & y[15];
  assign P[3][16] = x[3] & y[16];
  assign P[3][17] = x[3] & y[17];
  assign P[3][18] = x[3] & y[18];
  assign P[3][19] = x[3] & y[19];
  assign P[3][20] = x[3] & y[20];
  assign P[3][21] = x[3] & y[21];
  assign P[3][22] = x[3] & y[22];
  assign P[3][23] = x[3] & y[23];
  assign P[3][24] = x[3] & y[24];
  assign P[3][25] = x[3] & y[25];
  assign P[3][26] = x[3] & y[26];
  assign P[3][27] = x[3] & y[27];
  assign P[3][28] = x[3] & y[28];
  assign P[3][29] = x[3] & y[29];
  assign P[3][30] = x[3] & y[30];
  assign P[3][31] = x[3] & y[31];
  assign P[4][0] = x[4] & y[0];
  assign P[4][1] = x[4] & y[1];
  assign P[4][2] = x[4] & y[2];
  assign P[4][3] = x[4] & y[3];
  assign P[4][4] = x[4] & y[4];
  assign P[4][5] = x[4] & y[5];
  assign P[4][6] = x[4] & y[6];
  assign P[4][7] = x[4] & y[7];
  assign P[4][8] = x[4] & y[8];
  assign P[4][9] = x[4] & y[9];
  assign P[4][10] = x[4] & y[10];
  assign P[4][11] = x[4] & y[11];
  assign P[4][12] = x[4] & y[12];
  assign P[4][13] = x[4] & y[13];
  assign P[4][14] = x[4] & y[14];
  assign P[4][15] = x[4] & y[15];
  assign P[4][16] = x[4] & y[16];
  assign P[4][17] = x[4] & y[17];
  assign P[4][18] = x[4] & y[18];
  assign P[4][19] = x[4] & y[19];
  assign P[4][20] = x[4] & y[20];
  assign P[4][21] = x[4] & y[21];
  assign P[4][22] = x[4] & y[22];
  assign P[4][23] = x[4] & y[23];
  assign P[4][24] = x[4] & y[24];
  assign P[4][25] = x[4] & y[25];
  assign P[4][26] = x[4] & y[26];
  assign P[4][27] = x[4] & y[27];
  assign P[4][28] = x[4] & y[28];
  assign P[4][29] = x[4] & y[29];
  assign P[4][30] = x[4] & y[30];
  assign P[4][31] = x[4] & y[31];
  assign P[5][0] = x[5] & y[0];
  assign P[5][1] = x[5] & y[1];
  assign P[5][2] = x[5] & y[2];
  assign P[5][3] = x[5] & y[3];
  assign P[5][4] = x[5] & y[4];
  assign P[5][5] = x[5] & y[5];
  assign P[5][6] = x[5] & y[6];
  assign P[5][7] = x[5] & y[7];
  assign P[5][8] = x[5] & y[8];
  assign P[5][9] = x[5] & y[9];
  assign P[5][10] = x[5] & y[10];
  assign P[5][11] = x[5] & y[11];
  assign P[5][12] = x[5] & y[12];
  assign P[5][13] = x[5] & y[13];
  assign P[5][14] = x[5] & y[14];
  assign P[5][15] = x[5] & y[15];
  assign P[5][16] = x[5] & y[16];
  assign P[5][17] = x[5] & y[17];
  assign P[5][18] = x[5] & y[18];
  assign P[5][19] = x[5] & y[19];
  assign P[5][20] = x[5] & y[20];
  assign P[5][21] = x[5] & y[21];
  assign P[5][22] = x[5] & y[22];
  assign P[5][23] = x[5] & y[23];
  assign P[5][24] = x[5] & y[24];
  assign P[5][25] = x[5] & y[25];
  assign P[5][26] = x[5] & y[26];
  assign P[5][27] = x[5] & y[27];
  assign P[5][28] = x[5] & y[28];
  assign P[5][29] = x[5] & y[29];
  assign P[5][30] = x[5] & y[30];
  assign P[5][31] = x[5] & y[31];
  assign P[6][0] = x[6] & y[0];
  assign P[6][1] = x[6] & y[1];
  assign P[6][2] = x[6] & y[2];
  assign P[6][3] = x[6] & y[3];
  assign P[6][4] = x[6] & y[4];
  assign P[6][5] = x[6] & y[5];
  assign P[6][6] = x[6] & y[6];
  assign P[6][7] = x[6] & y[7];
  assign P[6][8] = x[6] & y[8];
  assign P[6][9] = x[6] & y[9];
  assign P[6][10] = x[6] & y[10];
  assign P[6][11] = x[6] & y[11];
  assign P[6][12] = x[6] & y[12];
  assign P[6][13] = x[6] & y[13];
  assign P[6][14] = x[6] & y[14];
  assign P[6][15] = x[6] & y[15];
  assign P[6][16] = x[6] & y[16];
  assign P[6][17] = x[6] & y[17];
  assign P[6][18] = x[6] & y[18];
  assign P[6][19] = x[6] & y[19];
  assign P[6][20] = x[6] & y[20];
  assign P[6][21] = x[6] & y[21];
  assign P[6][22] = x[6] & y[22];
  assign P[6][23] = x[6] & y[23];
  assign P[6][24] = x[6] & y[24];
  assign P[6][25] = x[6] & y[25];
  assign P[6][26] = x[6] & y[26];
  assign P[6][27] = x[6] & y[27];
  assign P[6][28] = x[6] & y[28];
  assign P[6][29] = x[6] & y[29];
  assign P[6][30] = x[6] & y[30];
  assign P[6][31] = x[6] & y[31];
  assign P[7][0] = x[7] & y[0];
  assign P[7][1] = x[7] & y[1];
  assign P[7][2] = x[7] & y[2];
  assign P[7][3] = x[7] & y[3];
  assign P[7][4] = x[7] & y[4];
  assign P[7][5] = x[7] & y[5];
  assign P[7][6] = x[7] & y[6];
  assign P[7][7] = x[7] & y[7];
  assign P[7][8] = x[7] & y[8];
  assign P[7][9] = x[7] & y[9];
  assign P[7][10] = x[7] & y[10];
  assign P[7][11] = x[7] & y[11];
  assign P[7][12] = x[7] & y[12];
  assign P[7][13] = x[7] & y[13];
  assign P[7][14] = x[7] & y[14];
  assign P[7][15] = x[7] & y[15];
  assign P[7][16] = x[7] & y[16];
  assign P[7][17] = x[7] & y[17];
  assign P[7][18] = x[7] & y[18];
  assign P[7][19] = x[7] & y[19];
  assign P[7][20] = x[7] & y[20];
  assign P[7][21] = x[7] & y[21];
  assign P[7][22] = x[7] & y[22];
  assign P[7][23] = x[7] & y[23];
  assign P[7][24] = x[7] & y[24];
  assign P[7][25] = x[7] & y[25];
  assign P[7][26] = x[7] & y[26];
  assign P[7][27] = x[7] & y[27];
  assign P[7][28] = x[7] & y[28];
  assign P[7][29] = x[7] & y[29];
  assign P[7][30] = x[7] & y[30];
  assign P[7][31] = x[7] & y[31];
  assign P[8][0] = x[8] & y[0];
  assign P[8][1] = x[8] & y[1];
  assign P[8][2] = x[8] & y[2];
  assign P[8][3] = x[8] & y[3];
  assign P[8][4] = x[8] & y[4];
  assign P[8][5] = x[8] & y[5];
  assign P[8][6] = x[8] & y[6];
  assign P[8][7] = x[8] & y[7];
  assign P[8][8] = x[8] & y[8];
  assign P[8][9] = x[8] & y[9];
  assign P[8][10] = x[8] & y[10];
  assign P[8][11] = x[8] & y[11];
  assign P[8][12] = x[8] & y[12];
  assign P[8][13] = x[8] & y[13];
  assign P[8][14] = x[8] & y[14];
  assign P[8][15] = x[8] & y[15];
  assign P[8][16] = x[8] & y[16];
  assign P[8][17] = x[8] & y[17];
  assign P[8][18] = x[8] & y[18];
  assign P[8][19] = x[8] & y[19];
  assign P[8][20] = x[8] & y[20];
  assign P[8][21] = x[8] & y[21];
  assign P[8][22] = x[8] & y[22];
  assign P[8][23] = x[8] & y[23];
  assign P[8][24] = x[8] & y[24];
  assign P[8][25] = x[8] & y[25];
  assign P[8][26] = x[8] & y[26];
  assign P[8][27] = x[8] & y[27];
  assign P[8][28] = x[8] & y[28];
  assign P[8][29] = x[8] & y[29];
  assign P[8][30] = x[8] & y[30];
  assign P[8][31] = x[8] & y[31];
  assign P[9][0] = x[9] & y[0];
  assign P[9][1] = x[9] & y[1];
  assign P[9][2] = x[9] & y[2];
  assign P[9][3] = x[9] & y[3];
  assign P[9][4] = x[9] & y[4];
  assign P[9][5] = x[9] & y[5];
  assign P[9][6] = x[9] & y[6];
  assign P[9][7] = x[9] & y[7];
  assign P[9][8] = x[9] & y[8];
  assign P[9][9] = x[9] & y[9];
  assign P[9][10] = x[9] & y[10];
  assign P[9][11] = x[9] & y[11];
  assign P[9][12] = x[9] & y[12];
  assign P[9][13] = x[9] & y[13];
  assign P[9][14] = x[9] & y[14];
  assign P[9][15] = x[9] & y[15];
  assign P[9][16] = x[9] & y[16];
  assign P[9][17] = x[9] & y[17];
  assign P[9][18] = x[9] & y[18];
  assign P[9][19] = x[9] & y[19];
  assign P[9][20] = x[9] & y[20];
  assign P[9][21] = x[9] & y[21];
  assign P[9][22] = x[9] & y[22];
  assign P[9][23] = x[9] & y[23];
  assign P[9][24] = x[9] & y[24];
  assign P[9][25] = x[9] & y[25];
  assign P[9][26] = x[9] & y[26];
  assign P[9][27] = x[9] & y[27];
  assign P[9][28] = x[9] & y[28];
  assign P[9][29] = x[9] & y[29];
  assign P[9][30] = x[9] & y[30];
  assign P[9][31] = x[9] & y[31];
  assign P[10][0] = x[10] & y[0];
  assign P[10][1] = x[10] & y[1];
  assign P[10][2] = x[10] & y[2];
  assign P[10][3] = x[10] & y[3];
  assign P[10][4] = x[10] & y[4];
  assign P[10][5] = x[10] & y[5];
  assign P[10][6] = x[10] & y[6];
  assign P[10][7] = x[10] & y[7];
  assign P[10][8] = x[10] & y[8];
  assign P[10][9] = x[10] & y[9];
  assign P[10][10] = x[10] & y[10];
  assign P[10][11] = x[10] & y[11];
  assign P[10][12] = x[10] & y[12];
  assign P[10][13] = x[10] & y[13];
  assign P[10][14] = x[10] & y[14];
  assign P[10][15] = x[10] & y[15];
  assign P[10][16] = x[10] & y[16];
  assign P[10][17] = x[10] & y[17];
  assign P[10][18] = x[10] & y[18];
  assign P[10][19] = x[10] & y[19];
  assign P[10][20] = x[10] & y[20];
  assign P[10][21] = x[10] & y[21];
  assign P[10][22] = x[10] & y[22];
  assign P[10][23] = x[10] & y[23];
  assign P[10][24] = x[10] & y[24];
  assign P[10][25] = x[10] & y[25];
  assign P[10][26] = x[10] & y[26];
  assign P[10][27] = x[10] & y[27];
  assign P[10][28] = x[10] & y[28];
  assign P[10][29] = x[10] & y[29];
  assign P[10][30] = x[10] & y[30];
  assign P[10][31] = x[10] & y[31];
  assign P[11][0] = x[11] & y[0];
  assign P[11][1] = x[11] & y[1];
  assign P[11][2] = x[11] & y[2];
  assign P[11][3] = x[11] & y[3];
  assign P[11][4] = x[11] & y[4];
  assign P[11][5] = x[11] & y[5];
  assign P[11][6] = x[11] & y[6];
  assign P[11][7] = x[11] & y[7];
  assign P[11][8] = x[11] & y[8];
  assign P[11][9] = x[11] & y[9];
  assign P[11][10] = x[11] & y[10];
  assign P[11][11] = x[11] & y[11];
  assign P[11][12] = x[11] & y[12];
  assign P[11][13] = x[11] & y[13];
  assign P[11][14] = x[11] & y[14];
  assign P[11][15] = x[11] & y[15];
  assign P[11][16] = x[11] & y[16];
  assign P[11][17] = x[11] & y[17];
  assign P[11][18] = x[11] & y[18];
  assign P[11][19] = x[11] & y[19];
  assign P[11][20] = x[11] & y[20];
  assign P[11][21] = x[11] & y[21];
  assign P[11][22] = x[11] & y[22];
  assign P[11][23] = x[11] & y[23];
  assign P[11][24] = x[11] & y[24];
  assign P[11][25] = x[11] & y[25];
  assign P[11][26] = x[11] & y[26];
  assign P[11][27] = x[11] & y[27];
  assign P[11][28] = x[11] & y[28];
  assign P[11][29] = x[11] & y[29];
  assign P[11][30] = x[11] & y[30];
  assign P[11][31] = x[11] & y[31];
  assign P[12][0] = x[12] & y[0];
  assign P[12][1] = x[12] & y[1];
  assign P[12][2] = x[12] & y[2];
  assign P[12][3] = x[12] & y[3];
  assign P[12][4] = x[12] & y[4];
  assign P[12][5] = x[12] & y[5];
  assign P[12][6] = x[12] & y[6];
  assign P[12][7] = x[12] & y[7];
  assign P[12][8] = x[12] & y[8];
  assign P[12][9] = x[12] & y[9];
  assign P[12][10] = x[12] & y[10];
  assign P[12][11] = x[12] & y[11];
  assign P[12][12] = x[12] & y[12];
  assign P[12][13] = x[12] & y[13];
  assign P[12][14] = x[12] & y[14];
  assign P[12][15] = x[12] & y[15];
  assign P[12][16] = x[12] & y[16];
  assign P[12][17] = x[12] & y[17];
  assign P[12][18] = x[12] & y[18];
  assign P[12][19] = x[12] & y[19];
  assign P[12][20] = x[12] & y[20];
  assign P[12][21] = x[12] & y[21];
  assign P[12][22] = x[12] & y[22];
  assign P[12][23] = x[12] & y[23];
  assign P[12][24] = x[12] & y[24];
  assign P[12][25] = x[12] & y[25];
  assign P[12][26] = x[12] & y[26];
  assign P[12][27] = x[12] & y[27];
  assign P[12][28] = x[12] & y[28];
  assign P[12][29] = x[12] & y[29];
  assign P[12][30] = x[12] & y[30];
  assign P[12][31] = x[12] & y[31];
  assign P[13][0] = x[13] & y[0];
  assign P[13][1] = x[13] & y[1];
  assign P[13][2] = x[13] & y[2];
  assign P[13][3] = x[13] & y[3];
  assign P[13][4] = x[13] & y[4];
  assign P[13][5] = x[13] & y[5];
  assign P[13][6] = x[13] & y[6];
  assign P[13][7] = x[13] & y[7];
  assign P[13][8] = x[13] & y[8];
  assign P[13][9] = x[13] & y[9];
  assign P[13][10] = x[13] & y[10];
  assign P[13][11] = x[13] & y[11];
  assign P[13][12] = x[13] & y[12];
  assign P[13][13] = x[13] & y[13];
  assign P[13][14] = x[13] & y[14];
  assign P[13][15] = x[13] & y[15];
  assign P[13][16] = x[13] & y[16];
  assign P[13][17] = x[13] & y[17];
  assign P[13][18] = x[13] & y[18];
  assign P[13][19] = x[13] & y[19];
  assign P[13][20] = x[13] & y[20];
  assign P[13][21] = x[13] & y[21];
  assign P[13][22] = x[13] & y[22];
  assign P[13][23] = x[13] & y[23];
  assign P[13][24] = x[13] & y[24];
  assign P[13][25] = x[13] & y[25];
  assign P[13][26] = x[13] & y[26];
  assign P[13][27] = x[13] & y[27];
  assign P[13][28] = x[13] & y[28];
  assign P[13][29] = x[13] & y[29];
  assign P[13][30] = x[13] & y[30];
  assign P[13][31] = x[13] & y[31];
  assign P[14][0] = x[14] & y[0];
  assign P[14][1] = x[14] & y[1];
  assign P[14][2] = x[14] & y[2];
  assign P[14][3] = x[14] & y[3];
  assign P[14][4] = x[14] & y[4];
  assign P[14][5] = x[14] & y[5];
  assign P[14][6] = x[14] & y[6];
  assign P[14][7] = x[14] & y[7];
  assign P[14][8] = x[14] & y[8];
  assign P[14][9] = x[14] & y[9];
  assign P[14][10] = x[14] & y[10];
  assign P[14][11] = x[14] & y[11];
  assign P[14][12] = x[14] & y[12];
  assign P[14][13] = x[14] & y[13];
  assign P[14][14] = x[14] & y[14];
  assign P[14][15] = x[14] & y[15];
  assign P[14][16] = x[14] & y[16];
  assign P[14][17] = x[14] & y[17];
  assign P[14][18] = x[14] & y[18];
  assign P[14][19] = x[14] & y[19];
  assign P[14][20] = x[14] & y[20];
  assign P[14][21] = x[14] & y[21];
  assign P[14][22] = x[14] & y[22];
  assign P[14][23] = x[14] & y[23];
  assign P[14][24] = x[14] & y[24];
  assign P[14][25] = x[14] & y[25];
  assign P[14][26] = x[14] & y[26];
  assign P[14][27] = x[14] & y[27];
  assign P[14][28] = x[14] & y[28];
  assign P[14][29] = x[14] & y[29];
  assign P[14][30] = x[14] & y[30];
  assign P[14][31] = x[14] & y[31];
  assign P[15][0] = x[15] & y[0];
  assign P[15][1] = x[15] & y[1];
  assign P[15][2] = x[15] & y[2];
  assign P[15][3] = x[15] & y[3];
  assign P[15][4] = x[15] & y[4];
  assign P[15][5] = x[15] & y[5];
  assign P[15][6] = x[15] & y[6];
  assign P[15][7] = x[15] & y[7];
  assign P[15][8] = x[15] & y[8];
  assign P[15][9] = x[15] & y[9];
  assign P[15][10] = x[15] & y[10];
  assign P[15][11] = x[15] & y[11];
  assign P[15][12] = x[15] & y[12];
  assign P[15][13] = x[15] & y[13];
  assign P[15][14] = x[15] & y[14];
  assign P[15][15] = x[15] & y[15];
  assign P[15][16] = x[15] & y[16];
  assign P[15][17] = x[15] & y[17];
  assign P[15][18] = x[15] & y[18];
  assign P[15][19] = x[15] & y[19];
  assign P[15][20] = x[15] & y[20];
  assign P[15][21] = x[15] & y[21];
  assign P[15][22] = x[15] & y[22];
  assign P[15][23] = x[15] & y[23];
  assign P[15][24] = x[15] & y[24];
  assign P[15][25] = x[15] & y[25];
  assign P[15][26] = x[15] & y[26];
  assign P[15][27] = x[15] & y[27];
  assign P[15][28] = x[15] & y[28];
  assign P[15][29] = x[15] & y[29];
  assign P[15][30] = x[15] & y[30];
  assign P[15][31] = x[15] & y[31];
  assign P[16][0] = x[16] & y[0];
  assign P[16][1] = x[16] & y[1];
  assign P[16][2] = x[16] & y[2];
  assign P[16][3] = x[16] & y[3];
  assign P[16][4] = x[16] & y[4];
  assign P[16][5] = x[16] & y[5];
  assign P[16][6] = x[16] & y[6];
  assign P[16][7] = x[16] & y[7];
  assign P[16][8] = x[16] & y[8];
  assign P[16][9] = x[16] & y[9];
  assign P[16][10] = x[16] & y[10];
  assign P[16][11] = x[16] & y[11];
  assign P[16][12] = x[16] & y[12];
  assign P[16][13] = x[16] & y[13];
  assign P[16][14] = x[16] & y[14];
  assign P[16][15] = x[16] & y[15];
  assign P[16][16] = x[16] & y[16];
  assign P[16][17] = x[16] & y[17];
  assign P[16][18] = x[16] & y[18];
  assign P[16][19] = x[16] & y[19];
  assign P[16][20] = x[16] & y[20];
  assign P[16][21] = x[16] & y[21];
  assign P[16][22] = x[16] & y[22];
  assign P[16][23] = x[16] & y[23];
  assign P[16][24] = x[16] & y[24];
  assign P[16][25] = x[16] & y[25];
  assign P[16][26] = x[16] & y[26];
  assign P[16][27] = x[16] & y[27];
  assign P[16][28] = x[16] & y[28];
  assign P[16][29] = x[16] & y[29];
  assign P[16][30] = x[16] & y[30];
  assign P[16][31] = x[16] & y[31];
  assign P[17][0] = x[17] & y[0];
  assign P[17][1] = x[17] & y[1];
  assign P[17][2] = x[17] & y[2];
  assign P[17][3] = x[17] & y[3];
  assign P[17][4] = x[17] & y[4];
  assign P[17][5] = x[17] & y[5];
  assign P[17][6] = x[17] & y[6];
  assign P[17][7] = x[17] & y[7];
  assign P[17][8] = x[17] & y[8];
  assign P[17][9] = x[17] & y[9];
  assign P[17][10] = x[17] & y[10];
  assign P[17][11] = x[17] & y[11];
  assign P[17][12] = x[17] & y[12];
  assign P[17][13] = x[17] & y[13];
  assign P[17][14] = x[17] & y[14];
  assign P[17][15] = x[17] & y[15];
  assign P[17][16] = x[17] & y[16];
  assign P[17][17] = x[17] & y[17];
  assign P[17][18] = x[17] & y[18];
  assign P[17][19] = x[17] & y[19];
  assign P[17][20] = x[17] & y[20];
  assign P[17][21] = x[17] & y[21];
  assign P[17][22] = x[17] & y[22];
  assign P[17][23] = x[17] & y[23];
  assign P[17][24] = x[17] & y[24];
  assign P[17][25] = x[17] & y[25];
  assign P[17][26] = x[17] & y[26];
  assign P[17][27] = x[17] & y[27];
  assign P[17][28] = x[17] & y[28];
  assign P[17][29] = x[17] & y[29];
  assign P[17][30] = x[17] & y[30];
  assign P[17][31] = x[17] & y[31];
  assign P[18][0] = x[18] & y[0];
  assign P[18][1] = x[18] & y[1];
  assign P[18][2] = x[18] & y[2];
  assign P[18][3] = x[18] & y[3];
  assign P[18][4] = x[18] & y[4];
  assign P[18][5] = x[18] & y[5];
  assign P[18][6] = x[18] & y[6];
  assign P[18][7] = x[18] & y[7];
  assign P[18][8] = x[18] & y[8];
  assign P[18][9] = x[18] & y[9];
  assign P[18][10] = x[18] & y[10];
  assign P[18][11] = x[18] & y[11];
  assign P[18][12] = x[18] & y[12];
  assign P[18][13] = x[18] & y[13];
  assign P[18][14] = x[18] & y[14];
  assign P[18][15] = x[18] & y[15];
  assign P[18][16] = x[18] & y[16];
  assign P[18][17] = x[18] & y[17];
  assign P[18][18] = x[18] & y[18];
  assign P[18][19] = x[18] & y[19];
  assign P[18][20] = x[18] & y[20];
  assign P[18][21] = x[18] & y[21];
  assign P[18][22] = x[18] & y[22];
  assign P[18][23] = x[18] & y[23];
  assign P[18][24] = x[18] & y[24];
  assign P[18][25] = x[18] & y[25];
  assign P[18][26] = x[18] & y[26];
  assign P[18][27] = x[18] & y[27];
  assign P[18][28] = x[18] & y[28];
  assign P[18][29] = x[18] & y[29];
  assign P[18][30] = x[18] & y[30];
  assign P[18][31] = x[18] & y[31];
  assign P[19][0] = x[19] & y[0];
  assign P[19][1] = x[19] & y[1];
  assign P[19][2] = x[19] & y[2];
  assign P[19][3] = x[19] & y[3];
  assign P[19][4] = x[19] & y[4];
  assign P[19][5] = x[19] & y[5];
  assign P[19][6] = x[19] & y[6];
  assign P[19][7] = x[19] & y[7];
  assign P[19][8] = x[19] & y[8];
  assign P[19][9] = x[19] & y[9];
  assign P[19][10] = x[19] & y[10];
  assign P[19][11] = x[19] & y[11];
  assign P[19][12] = x[19] & y[12];
  assign P[19][13] = x[19] & y[13];
  assign P[19][14] = x[19] & y[14];
  assign P[19][15] = x[19] & y[15];
  assign P[19][16] = x[19] & y[16];
  assign P[19][17] = x[19] & y[17];
  assign P[19][18] = x[19] & y[18];
  assign P[19][19] = x[19] & y[19];
  assign P[19][20] = x[19] & y[20];
  assign P[19][21] = x[19] & y[21];
  assign P[19][22] = x[19] & y[22];
  assign P[19][23] = x[19] & y[23];
  assign P[19][24] = x[19] & y[24];
  assign P[19][25] = x[19] & y[25];
  assign P[19][26] = x[19] & y[26];
  assign P[19][27] = x[19] & y[27];
  assign P[19][28] = x[19] & y[28];
  assign P[19][29] = x[19] & y[29];
  assign P[19][30] = x[19] & y[30];
  assign P[19][31] = x[19] & y[31];
  assign P[20][0] = x[20] & y[0];
  assign P[20][1] = x[20] & y[1];
  assign P[20][2] = x[20] & y[2];
  assign P[20][3] = x[20] & y[3];
  assign P[20][4] = x[20] & y[4];
  assign P[20][5] = x[20] & y[5];
  assign P[20][6] = x[20] & y[6];
  assign P[20][7] = x[20] & y[7];
  assign P[20][8] = x[20] & y[8];
  assign P[20][9] = x[20] & y[9];
  assign P[20][10] = x[20] & y[10];
  assign P[20][11] = x[20] & y[11];
  assign P[20][12] = x[20] & y[12];
  assign P[20][13] = x[20] & y[13];
  assign P[20][14] = x[20] & y[14];
  assign P[20][15] = x[20] & y[15];
  assign P[20][16] = x[20] & y[16];
  assign P[20][17] = x[20] & y[17];
  assign P[20][18] = x[20] & y[18];
  assign P[20][19] = x[20] & y[19];
  assign P[20][20] = x[20] & y[20];
  assign P[20][21] = x[20] & y[21];
  assign P[20][22] = x[20] & y[22];
  assign P[20][23] = x[20] & y[23];
  assign P[20][24] = x[20] & y[24];
  assign P[20][25] = x[20] & y[25];
  assign P[20][26] = x[20] & y[26];
  assign P[20][27] = x[20] & y[27];
  assign P[20][28] = x[20] & y[28];
  assign P[20][29] = x[20] & y[29];
  assign P[20][30] = x[20] & y[30];
  assign P[20][31] = x[20] & y[31];
  assign P[21][0] = x[21] & y[0];
  assign P[21][1] = x[21] & y[1];
  assign P[21][2] = x[21] & y[2];
  assign P[21][3] = x[21] & y[3];
  assign P[21][4] = x[21] & y[4];
  assign P[21][5] = x[21] & y[5];
  assign P[21][6] = x[21] & y[6];
  assign P[21][7] = x[21] & y[7];
  assign P[21][8] = x[21] & y[8];
  assign P[21][9] = x[21] & y[9];
  assign P[21][10] = x[21] & y[10];
  assign P[21][11] = x[21] & y[11];
  assign P[21][12] = x[21] & y[12];
  assign P[21][13] = x[21] & y[13];
  assign P[21][14] = x[21] & y[14];
  assign P[21][15] = x[21] & y[15];
  assign P[21][16] = x[21] & y[16];
  assign P[21][17] = x[21] & y[17];
  assign P[21][18] = x[21] & y[18];
  assign P[21][19] = x[21] & y[19];
  assign P[21][20] = x[21] & y[20];
  assign P[21][21] = x[21] & y[21];
  assign P[21][22] = x[21] & y[22];
  assign P[21][23] = x[21] & y[23];
  assign P[21][24] = x[21] & y[24];
  assign P[21][25] = x[21] & y[25];
  assign P[21][26] = x[21] & y[26];
  assign P[21][27] = x[21] & y[27];
  assign P[21][28] = x[21] & y[28];
  assign P[21][29] = x[21] & y[29];
  assign P[21][30] = x[21] & y[30];
  assign P[21][31] = x[21] & y[31];
  assign P[22][0] = x[22] & y[0];
  assign P[22][1] = x[22] & y[1];
  assign P[22][2] = x[22] & y[2];
  assign P[22][3] = x[22] & y[3];
  assign P[22][4] = x[22] & y[4];
  assign P[22][5] = x[22] & y[5];
  assign P[22][6] = x[22] & y[6];
  assign P[22][7] = x[22] & y[7];
  assign P[22][8] = x[22] & y[8];
  assign P[22][9] = x[22] & y[9];
  assign P[22][10] = x[22] & y[10];
  assign P[22][11] = x[22] & y[11];
  assign P[22][12] = x[22] & y[12];
  assign P[22][13] = x[22] & y[13];
  assign P[22][14] = x[22] & y[14];
  assign P[22][15] = x[22] & y[15];
  assign P[22][16] = x[22] & y[16];
  assign P[22][17] = x[22] & y[17];
  assign P[22][18] = x[22] & y[18];
  assign P[22][19] = x[22] & y[19];
  assign P[22][20] = x[22] & y[20];
  assign P[22][21] = x[22] & y[21];
  assign P[22][22] = x[22] & y[22];
  assign P[22][23] = x[22] & y[23];
  assign P[22][24] = x[22] & y[24];
  assign P[22][25] = x[22] & y[25];
  assign P[22][26] = x[22] & y[26];
  assign P[22][27] = x[22] & y[27];
  assign P[22][28] = x[22] & y[28];
  assign P[22][29] = x[22] & y[29];
  assign P[22][30] = x[22] & y[30];
  assign P[22][31] = x[22] & y[31];
  assign P[23][0] = x[23] & y[0];
  assign P[23][1] = x[23] & y[1];
  assign P[23][2] = x[23] & y[2];
  assign P[23][3] = x[23] & y[3];
  assign P[23][4] = x[23] & y[4];
  assign P[23][5] = x[23] & y[5];
  assign P[23][6] = x[23] & y[6];
  assign P[23][7] = x[23] & y[7];
  assign P[23][8] = x[23] & y[8];
  assign P[23][9] = x[23] & y[9];
  assign P[23][10] = x[23] & y[10];
  assign P[23][11] = x[23] & y[11];
  assign P[23][12] = x[23] & y[12];
  assign P[23][13] = x[23] & y[13];
  assign P[23][14] = x[23] & y[14];
  assign P[23][15] = x[23] & y[15];
  assign P[23][16] = x[23] & y[16];
  assign P[23][17] = x[23] & y[17];
  assign P[23][18] = x[23] & y[18];
  assign P[23][19] = x[23] & y[19];
  assign P[23][20] = x[23] & y[20];
  assign P[23][21] = x[23] & y[21];
  assign P[23][22] = x[23] & y[22];
  assign P[23][23] = x[23] & y[23];
  assign P[23][24] = x[23] & y[24];
  assign P[23][25] = x[23] & y[25];
  assign P[23][26] = x[23] & y[26];
  assign P[23][27] = x[23] & y[27];
  assign P[23][28] = x[23] & y[28];
  assign P[23][29] = x[23] & y[29];
  assign P[23][30] = x[23] & y[30];
  assign P[23][31] = x[23] & y[31];
  assign P[24][0] = x[24] & y[0];
  assign P[24][1] = x[24] & y[1];
  assign P[24][2] = x[24] & y[2];
  assign P[24][3] = x[24] & y[3];
  assign P[24][4] = x[24] & y[4];
  assign P[24][5] = x[24] & y[5];
  assign P[24][6] = x[24] & y[6];
  assign P[24][7] = x[24] & y[7];
  assign P[24][8] = x[24] & y[8];
  assign P[24][9] = x[24] & y[9];
  assign P[24][10] = x[24] & y[10];
  assign P[24][11] = x[24] & y[11];
  assign P[24][12] = x[24] & y[12];
  assign P[24][13] = x[24] & y[13];
  assign P[24][14] = x[24] & y[14];
  assign P[24][15] = x[24] & y[15];
  assign P[24][16] = x[24] & y[16];
  assign P[24][17] = x[24] & y[17];
  assign P[24][18] = x[24] & y[18];
  assign P[24][19] = x[24] & y[19];
  assign P[24][20] = x[24] & y[20];
  assign P[24][21] = x[24] & y[21];
  assign P[24][22] = x[24] & y[22];
  assign P[24][23] = x[24] & y[23];
  assign P[24][24] = x[24] & y[24];
  assign P[24][25] = x[24] & y[25];
  assign P[24][26] = x[24] & y[26];
  assign P[24][27] = x[24] & y[27];
  assign P[24][28] = x[24] & y[28];
  assign P[24][29] = x[24] & y[29];
  assign P[24][30] = x[24] & y[30];
  assign P[24][31] = x[24] & y[31];
  assign P[25][0] = x[25] & y[0];
  assign P[25][1] = x[25] & y[1];
  assign P[25][2] = x[25] & y[2];
  assign P[25][3] = x[25] & y[3];
  assign P[25][4] = x[25] & y[4];
  assign P[25][5] = x[25] & y[5];
  assign P[25][6] = x[25] & y[6];
  assign P[25][7] = x[25] & y[7];
  assign P[25][8] = x[25] & y[8];
  assign P[25][9] = x[25] & y[9];
  assign P[25][10] = x[25] & y[10];
  assign P[25][11] = x[25] & y[11];
  assign P[25][12] = x[25] & y[12];
  assign P[25][13] = x[25] & y[13];
  assign P[25][14] = x[25] & y[14];
  assign P[25][15] = x[25] & y[15];
  assign P[25][16] = x[25] & y[16];
  assign P[25][17] = x[25] & y[17];
  assign P[25][18] = x[25] & y[18];
  assign P[25][19] = x[25] & y[19];
  assign P[25][20] = x[25] & y[20];
  assign P[25][21] = x[25] & y[21];
  assign P[25][22] = x[25] & y[22];
  assign P[25][23] = x[25] & y[23];
  assign P[25][24] = x[25] & y[24];
  assign P[25][25] = x[25] & y[25];
  assign P[25][26] = x[25] & y[26];
  assign P[25][27] = x[25] & y[27];
  assign P[25][28] = x[25] & y[28];
  assign P[25][29] = x[25] & y[29];
  assign P[25][30] = x[25] & y[30];
  assign P[25][31] = x[25] & y[31];
  assign P[26][0] = x[26] & y[0];
  assign P[26][1] = x[26] & y[1];
  assign P[26][2] = x[26] & y[2];
  assign P[26][3] = x[26] & y[3];
  assign P[26][4] = x[26] & y[4];
  assign P[26][5] = x[26] & y[5];
  assign P[26][6] = x[26] & y[6];
  assign P[26][7] = x[26] & y[7];
  assign P[26][8] = x[26] & y[8];
  assign P[26][9] = x[26] & y[9];
  assign P[26][10] = x[26] & y[10];
  assign P[26][11] = x[26] & y[11];
  assign P[26][12] = x[26] & y[12];
  assign P[26][13] = x[26] & y[13];
  assign P[26][14] = x[26] & y[14];
  assign P[26][15] = x[26] & y[15];
  assign P[26][16] = x[26] & y[16];
  assign P[26][17] = x[26] & y[17];
  assign P[26][18] = x[26] & y[18];
  assign P[26][19] = x[26] & y[19];
  assign P[26][20] = x[26] & y[20];
  assign P[26][21] = x[26] & y[21];
  assign P[26][22] = x[26] & y[22];
  assign P[26][23] = x[26] & y[23];
  assign P[26][24] = x[26] & y[24];
  assign P[26][25] = x[26] & y[25];
  assign P[26][26] = x[26] & y[26];
  assign P[26][27] = x[26] & y[27];
  assign P[26][28] = x[26] & y[28];
  assign P[26][29] = x[26] & y[29];
  assign P[26][30] = x[26] & y[30];
  assign P[26][31] = x[26] & y[31];
  assign P[27][0] = x[27] & y[0];
  assign P[27][1] = x[27] & y[1];
  assign P[27][2] = x[27] & y[2];
  assign P[27][3] = x[27] & y[3];
  assign P[27][4] = x[27] & y[4];
  assign P[27][5] = x[27] & y[5];
  assign P[27][6] = x[27] & y[6];
  assign P[27][7] = x[27] & y[7];
  assign P[27][8] = x[27] & y[8];
  assign P[27][9] = x[27] & y[9];
  assign P[27][10] = x[27] & y[10];
  assign P[27][11] = x[27] & y[11];
  assign P[27][12] = x[27] & y[12];
  assign P[27][13] = x[27] & y[13];
  assign P[27][14] = x[27] & y[14];
  assign P[27][15] = x[27] & y[15];
  assign P[27][16] = x[27] & y[16];
  assign P[27][17] = x[27] & y[17];
  assign P[27][18] = x[27] & y[18];
  assign P[27][19] = x[27] & y[19];
  assign P[27][20] = x[27] & y[20];
  assign P[27][21] = x[27] & y[21];
  assign P[27][22] = x[27] & y[22];
  assign P[27][23] = x[27] & y[23];
  assign P[27][24] = x[27] & y[24];
  assign P[27][25] = x[27] & y[25];
  assign P[27][26] = x[27] & y[26];
  assign P[27][27] = x[27] & y[27];
  assign P[27][28] = x[27] & y[28];
  assign P[27][29] = x[27] & y[29];
  assign P[27][30] = x[27] & y[30];
  assign P[27][31] = x[27] & y[31];
  assign P[28][0] = x[28] & y[0];
  assign P[28][1] = x[28] & y[1];
  assign P[28][2] = x[28] & y[2];
  assign P[28][3] = x[28] & y[3];
  assign P[28][4] = x[28] & y[4];
  assign P[28][5] = x[28] & y[5];
  assign P[28][6] = x[28] & y[6];
  assign P[28][7] = x[28] & y[7];
  assign P[28][8] = x[28] & y[8];
  assign P[28][9] = x[28] & y[9];
  assign P[28][10] = x[28] & y[10];
  assign P[28][11] = x[28] & y[11];
  assign P[28][12] = x[28] & y[12];
  assign P[28][13] = x[28] & y[13];
  assign P[28][14] = x[28] & y[14];
  assign P[28][15] = x[28] & y[15];
  assign P[28][16] = x[28] & y[16];
  assign P[28][17] = x[28] & y[17];
  assign P[28][18] = x[28] & y[18];
  assign P[28][19] = x[28] & y[19];
  assign P[28][20] = x[28] & y[20];
  assign P[28][21] = x[28] & y[21];
  assign P[28][22] = x[28] & y[22];
  assign P[28][23] = x[28] & y[23];
  assign P[28][24] = x[28] & y[24];
  assign P[28][25] = x[28] & y[25];
  assign P[28][26] = x[28] & y[26];
  assign P[28][27] = x[28] & y[27];
  assign P[28][28] = x[28] & y[28];
  assign P[28][29] = x[28] & y[29];
  assign P[28][30] = x[28] & y[30];
  assign P[28][31] = x[28] & y[31];
  assign P[29][0] = x[29] & y[0];
  assign P[29][1] = x[29] & y[1];
  assign P[29][2] = x[29] & y[2];
  assign P[29][3] = x[29] & y[3];
  assign P[29][4] = x[29] & y[4];
  assign P[29][5] = x[29] & y[5];
  assign P[29][6] = x[29] & y[6];
  assign P[29][7] = x[29] & y[7];
  assign P[29][8] = x[29] & y[8];
  assign P[29][9] = x[29] & y[9];
  assign P[29][10] = x[29] & y[10];
  assign P[29][11] = x[29] & y[11];
  assign P[29][12] = x[29] & y[12];
  assign P[29][13] = x[29] & y[13];
  assign P[29][14] = x[29] & y[14];
  assign P[29][15] = x[29] & y[15];
  assign P[29][16] = x[29] & y[16];
  assign P[29][17] = x[29] & y[17];
  assign P[29][18] = x[29] & y[18];
  assign P[29][19] = x[29] & y[19];
  assign P[29][20] = x[29] & y[20];
  assign P[29][21] = x[29] & y[21];
  assign P[29][22] = x[29] & y[22];
  assign P[29][23] = x[29] & y[23];
  assign P[29][24] = x[29] & y[24];
  assign P[29][25] = x[29] & y[25];
  assign P[29][26] = x[29] & y[26];
  assign P[29][27] = x[29] & y[27];
  assign P[29][28] = x[29] & y[28];
  assign P[29][29] = x[29] & y[29];
  assign P[29][30] = x[29] & y[30];
  assign P[29][31] = x[29] & y[31];
  assign P[30][0] = x[30] & y[0];
  assign P[30][1] = x[30] & y[1];
  assign P[30][2] = x[30] & y[2];
  assign P[30][3] = x[30] & y[3];
  assign P[30][4] = x[30] & y[4];
  assign P[30][5] = x[30] & y[5];
  assign P[30][6] = x[30] & y[6];
  assign P[30][7] = x[30] & y[7];
  assign P[30][8] = x[30] & y[8];
  assign P[30][9] = x[30] & y[9];
  assign P[30][10] = x[30] & y[10];
  assign P[30][11] = x[30] & y[11];
  assign P[30][12] = x[30] & y[12];
  assign P[30][13] = x[30] & y[13];
  assign P[30][14] = x[30] & y[14];
  assign P[30][15] = x[30] & y[15];
  assign P[30][16] = x[30] & y[16];
  assign P[30][17] = x[30] & y[17];
  assign P[30][18] = x[30] & y[18];
  assign P[30][19] = x[30] & y[19];
  assign P[30][20] = x[30] & y[20];
  assign P[30][21] = x[30] & y[21];
  assign P[30][22] = x[30] & y[22];
  assign P[30][23] = x[30] & y[23];
  assign P[30][24] = x[30] & y[24];
  assign P[30][25] = x[30] & y[25];
  assign P[30][26] = x[30] & y[26];
  assign P[30][27] = x[30] & y[27];
  assign P[30][28] = x[30] & y[28];
  assign P[30][29] = x[30] & y[29];
  assign P[30][30] = x[30] & y[30];
  assign P[30][31] = x[30] & y[31];
  assign P[31][0] = x[31] & y[0];
  assign P[31][1] = x[31] & y[1];
  assign P[31][2] = x[31] & y[2];
  assign P[31][3] = x[31] & y[3];
  assign P[31][4] = x[31] & y[4];
  assign P[31][5] = x[31] & y[5];
  assign P[31][6] = x[31] & y[6];
  assign P[31][7] = x[31] & y[7];
  assign P[31][8] = x[31] & y[8];
  assign P[31][9] = x[31] & y[9];
  assign P[31][10] = x[31] & y[10];
  assign P[31][11] = x[31] & y[11];
  assign P[31][12] = x[31] & y[12];
  assign P[31][13] = x[31] & y[13];
  assign P[31][14] = x[31] & y[14];
  assign P[31][15] = x[31] & y[15];
  assign P[31][16] = x[31] & y[16];
  assign P[31][17] = x[31] & y[17];
  assign P[31][18] = x[31] & y[18];
  assign P[31][19] = x[31] & y[19];
  assign P[31][20] = x[31] & y[20];
  assign P[31][21] = x[31] & y[21];
  assign P[31][22] = x[31] & y[22];
  assign P[31][23] = x[31] & y[23];
  assign P[31][24] = x[31] & y[24];
  assign P[31][25] = x[31] & y[25];
  assign P[31][26] = x[31] & y[26];
  assign P[31][27] = x[31] & y[27];
  assign P[31][28] = x[31] & y[28];
  assign P[31][29] = x[31] & y[29];
  assign P[31][30] = x[31] & y[30];
  assign P[31][31] = x[31] & y[31];

  ha HA_00000000 (P[0][28],P[1][27],S[0],C[0]);
  fa FA_00000001 (P[0][29],P[1][28],P[2][27],S[1],C[1]);
  ha HA_00000002 (P[3][26],P[4][25],S[2],C[2]);
  fa FA_00000003 (P[0][30],P[1][29],P[2][28],S[3],C[3]);
  fa FA_00000004 (P[3][27],P[4][26],P[5][25],S[4],C[4]);
  ha HA_00000005 (P[6][24],P[7][23],S[5],C[5]);
  fa FA_00000006 (P[0][31],P[1][30],P[2][29],S[6],C[6]);
  fa FA_00000007 (P[3][28],P[4][27],P[5][26],S[7],C[7]);
  fa FA_00000008 (P[6][25],P[7][24],P[8][23],S[8],C[8]);
  ha HA_00000009 (P[9][22],P[10][21],S[9],C[9]);
  fa FA_00000010 (P[1][31],P[2][30],P[3][29],S[10],C[10]);
  fa FA_00000011 (P[4][28],P[5][27],P[6][26],S[11],C[11]);
  fa FA_00000012 (P[7][25],P[8][24],P[9][23],S[12],C[12]);
  ha HA_00000013 (P[10][22],P[11][21],S[13],C[13]);
  fa FA_00000014 (P[2][31],P[3][30],P[4][29],S[14],C[14]);
  fa FA_00000015 (P[5][28],P[6][27],P[7][26],S[15],C[15]);
  fa FA_00000016 (P[8][25],P[9][24],P[10][23],S[16],C[16]);
  fa FA_00000017 (P[3][31],P[4][30],P[5][29],S[17],C[17]);
  fa FA_00000018 (P[6][28],P[7][27],P[8][26],S[18],C[18]);
  fa FA_00000019 (P[4][31],P[5][30],P[6][29],S[19],C[19]);
  ha HA_00000020 (P[0][19],P[1][18],S[20],C[20]);
  fa FA_00000021 (P[0][20],P[1][19],P[2][18],S[21],C[21]);
  ha HA_00000022 (P[3][17],P[4][16],S[22],C[22]);
  fa FA_00000023 (P[0][21],P[1][20],P[2][19],S[23],C[23]);
  fa FA_00000024 (P[3][18],P[4][17],P[5][16],S[24],C[24]);
  ha HA_00000025 (P[6][15],P[7][14],S[25],C[25]);
  fa FA_00000026 (P[0][22],P[1][21],P[2][20],S[26],C[26]);
  fa FA_00000027 (P[3][19],P[4][18],P[5][17],S[27],C[27]);
  fa FA_00000028 (P[6][16],P[7][15],P[8][14],S[28],C[28]);
  ha HA_00000029 (P[9][13],P[10][12],S[29],C[29]);
  fa FA_00000030 (P[0][23],P[1][22],P[2][21],S[30],C[30]);
  fa FA_00000031 (P[3][20],P[4][19],P[5][18],S[31],C[31]);
  fa FA_00000032 (P[6][17],P[7][16],P[8][15],S[32],C[32]);
  fa FA_00000033 (P[9][14],P[10][13],P[11][12],S[33],C[33]);
  ha HA_00000034 (P[12][11],P[13][10],S[34],C[34]);
  fa FA_00000035 (P[0][24],P[1][23],P[2][22],S[35],C[35]);
  fa FA_00000036 (P[3][21],P[4][20],P[5][19],S[36],C[36]);
  fa FA_00000037 (P[6][18],P[7][17],P[8][16],S[37],C[37]);
  fa FA_00000038 (P[9][15],P[10][14],P[11][13],S[38],C[38]);
  fa FA_00000039 (P[12][12],P[13][11],P[14][10],S[39],C[39]);
  ha HA_00000040 (P[15][9],P[16][8],S[40],C[40]);
  fa FA_00000041 (P[0][25],P[1][24],P[2][23],S[41],C[41]);
  fa FA_00000042 (P[3][22],P[4][21],P[5][20],S[42],C[42]);
  fa FA_00000043 (P[6][19],P[7][18],P[8][17],S[43],C[43]);
  fa FA_00000044 (P[9][16],P[10][15],P[11][14],S[44],C[44]);
  fa FA_00000045 (P[12][13],P[13][12],P[14][11],S[45],C[45]);
  fa FA_00000046 (P[15][10],P[16][9],P[17][8],S[46],C[46]);
  ha HA_00000047 (P[18][7],P[19][6],S[47],C[47]);
  fa FA_00000048 (P[0][26],P[1][25],P[2][24],S[48],C[48]);
  fa FA_00000049 (P[3][23],P[4][22],P[5][21],S[49],C[49]);
  fa FA_00000050 (P[6][20],P[7][19],P[8][18],S[50],C[50]);
  fa FA_00000051 (P[9][17],P[10][16],P[11][15],S[51],C[51]);
  fa FA_00000052 (P[12][14],P[13][13],P[14][12],S[52],C[52]);
  fa FA_00000053 (P[15][11],P[16][10],P[17][9],S[53],C[53]);
  fa FA_00000054 (P[18][8],P[19][7],P[20][6],S[54],C[54]);
  ha HA_00000055 (P[21][5],P[22][4],S[55],C[55]);
  fa FA_00000056 (P[0][27],P[1][26],P[2][25],S[56],C[56]);
  fa FA_00000057 (P[3][24],P[4][23],P[5][22],S[57],C[57]);
  fa FA_00000058 (P[6][21],P[7][20],P[8][19],S[58],C[58]);
  fa FA_00000059 (P[9][18],P[10][17],P[11][16],S[59],C[59]);
  fa FA_00000060 (P[12][15],P[13][14],P[14][13],S[60],C[60]);
  fa FA_00000061 (P[15][12],P[16][11],P[17][10],S[61],C[61]);
  fa FA_00000062 (P[18][9],P[19][8],P[20][7],S[62],C[62]);
  fa FA_00000063 (P[21][6],P[22][5],P[23][4],S[63],C[63]);
  ha HA_00000064 (P[24][3],P[25][2],S[64],C[64]);
  fa FA_00000065 (S[0],P[2][26],P[3][25],S[65],C[65]);
  fa FA_00000066 (P[4][24],P[5][23],P[6][22],S[66],C[66]);
  fa FA_00000067 (P[7][21],P[8][20],P[9][19],S[67],C[67]);
  fa FA_00000068 (P[10][18],P[11][17],P[12][16],S[68],C[68]);
  fa FA_00000069 (P[13][15],P[14][14],P[15][13],S[69],C[69]);
  fa FA_00000070 (P[16][12],P[17][11],P[18][10],S[70],C[70]);
  fa FA_00000071 (P[19][9],P[20][8],P[21][7],S[71],C[71]);
  fa FA_00000072 (P[22][6],P[23][5],P[24][4],S[72],C[72]);
  fa FA_00000073 (P[25][3],P[26][2],P[27][1],S[73],C[73]);
  fa FA_00000074 (S[1],C[0],S[2],S[74],C[74]);
  fa FA_00000075 (P[5][24],P[6][23],P[7][22],S[75],C[75]);
  fa FA_00000076 (P[8][21],P[9][20],P[10][19],S[76],C[76]);
  fa FA_00000077 (P[11][18],P[12][17],P[13][16],S[77],C[77]);
  fa FA_00000078 (P[14][15],P[15][14],P[16][13],S[78],C[78]);
  fa FA_00000079 (P[17][12],P[18][11],P[19][10],S[79],C[79]);
  fa FA_00000080 (P[20][9],P[21][8],P[22][7],S[80],C[80]);
  fa FA_00000081 (P[23][6],P[24][5],P[25][4],S[81],C[81]);
  fa FA_00000082 (P[26][3],P[27][2],P[28][1],S[82],C[82]);
  fa FA_00000083 (S[3],C[1],S[4],S[83],C[83]);
  fa FA_00000084 (C[2],S[5],P[8][22],S[84],C[84]);
  fa FA_00000085 (P[9][21],P[10][20],P[11][19],S[85],C[85]);
  fa FA_00000086 (P[12][18],P[13][17],P[14][16],S[86],C[86]);
  fa FA_00000087 (P[15][15],P[16][14],P[17][13],S[87],C[87]);
  fa FA_00000088 (P[18][12],P[19][11],P[20][10],S[88],C[88]);
  fa FA_00000089 (P[21][9],P[22][8],P[23][7],S[89],C[89]);
  fa FA_00000090 (P[24][6],P[25][5],P[26][4],S[90],C[90]);
  fa FA_00000091 (P[27][3],P[28][2],P[29][1],S[91],C[91]);
  fa FA_00000092 (S[6],C[3],S[7],S[92],C[92]);
  fa FA_00000093 (C[4],S[8],C[5],S[93],C[93]);
  fa FA_00000094 (S[9],P[11][20],P[12][19],S[94],C[94]);
  fa FA_00000095 (P[13][18],P[14][17],P[15][16],S[95],C[95]);
  fa FA_00000096 (P[16][15],P[17][14],P[18][13],S[96],C[96]);
  fa FA_00000097 (P[19][12],P[20][11],P[21][10],S[97],C[97]);
  fa FA_00000098 (P[22][9],P[23][8],P[24][7],S[98],C[98]);
  fa FA_00000099 (P[25][6],P[26][5],P[27][4],S[99],C[99]);
  fa FA_00000100 (P[28][3],P[29][2],P[30][1],S[100],C[100]);
  fa FA_00000101 (S[10],C[6],S[11],S[101],C[101]);
  fa FA_00000102 (C[7],S[12],C[8],S[102],C[102]);
  fa FA_00000103 (S[13],C[9],P[12][20],S[103],C[103]);
  fa FA_00000104 (P[13][19],P[14][18],P[15][17],S[104],C[104]);
  fa FA_00000105 (P[16][16],P[17][15],P[18][14],S[105],C[105]);
  fa FA_00000106 (P[19][13],P[20][12],P[21][11],S[106],C[106]);
  fa FA_00000107 (P[22][10],P[23][9],P[24][8],S[107],C[107]);
  fa FA_00000108 (P[25][7],P[26][6],P[27][5],S[108],C[108]);
  fa FA_00000109 (P[28][4],P[29][3],P[30][2],S[109],C[109]);
  fa FA_00000110 (S[14],C[10],S[15],S[110],C[110]);
  fa FA_00000111 (C[11],S[16],C[12],S[111],C[111]);
  fa FA_00000112 (C[13],P[11][22],P[12][21],S[112],C[112]);
  fa FA_00000113 (P[13][20],P[14][19],P[15][18],S[113],C[113]);
  fa FA_00000114 (P[16][17],P[17][16],P[18][15],S[114],C[114]);
  fa FA_00000115 (P[19][14],P[20][13],P[21][12],S[115],C[115]);
  fa FA_00000116 (P[22][11],P[23][10],P[24][9],S[116],C[116]);
  fa FA_00000117 (P[25][8],P[26][7],P[27][6],S[117],C[117]);
  fa FA_00000118 (P[28][5],P[29][4],P[30][3],S[118],C[118]);
  fa FA_00000119 (S[17],C[14],S[18],S[119],C[119]);
  fa FA_00000120 (C[15],C[16],P[9][25],S[120],C[120]);
  fa FA_00000121 (P[10][24],P[11][23],P[12][22],S[121],C[121]);
  fa FA_00000122 (P[13][21],P[14][20],P[15][19],S[122],C[122]);
  fa FA_00000123 (P[16][18],P[17][17],P[18][16],S[123],C[123]);
  fa FA_00000124 (P[19][15],P[20][14],P[21][13],S[124],C[124]);
  fa FA_00000125 (P[22][12],P[23][11],P[24][10],S[125],C[125]);
  fa FA_00000126 (P[25][9],P[26][8],P[27][7],S[126],C[126]);
  fa FA_00000127 (P[28][6],P[29][5],P[30][4],S[127],C[127]);
  fa FA_00000128 (S[19],C[17],C[18],S[128],C[128]);
  fa FA_00000129 (P[7][28],P[8][27],P[9][26],S[129],C[129]);
  fa FA_00000130 (P[10][25],P[11][24],P[12][23],S[130],C[130]);
  fa FA_00000131 (P[13][22],P[14][21],P[15][20],S[131],C[131]);
  fa FA_00000132 (P[16][19],P[17][18],P[18][17],S[132],C[132]);
  fa FA_00000133 (P[19][16],P[20][15],P[21][14],S[133],C[133]);
  fa FA_00000134 (P[22][13],P[23][12],P[24][11],S[134],C[134]);
  fa FA_00000135 (P[25][10],P[26][9],P[27][8],S[135],C[135]);
  fa FA_00000136 (P[28][7],P[29][6],P[30][5],S[136],C[136]);
  fa FA_00000137 (C[19],P[5][31],P[6][30],S[137],C[137]);
  fa FA_00000138 (P[7][29],P[8][28],P[9][27],S[138],C[138]);
  fa FA_00000139 (P[10][26],P[11][25],P[12][24],S[139],C[139]);
  fa FA_00000140 (P[13][23],P[14][22],P[15][21],S[140],C[140]);
  fa FA_00000141 (P[16][20],P[17][19],P[18][18],S[141],C[141]);
  fa FA_00000142 (P[19][17],P[20][16],P[21][15],S[142],C[142]);
  fa FA_00000143 (P[22][14],P[23][13],P[24][12],S[143],C[143]);
  fa FA_00000144 (P[25][11],P[26][10],P[27][9],S[144],C[144]);
  fa FA_00000145 (P[28][8],P[29][7],P[30][6],S[145],C[145]);
  fa FA_00000146 (P[6][31],P[7][30],P[8][29],S[146],C[146]);
  fa FA_00000147 (P[9][28],P[10][27],P[11][26],S[147],C[147]);
  fa FA_00000148 (P[12][25],P[13][24],P[14][23],S[148],C[148]);
  fa FA_00000149 (P[15][22],P[16][21],P[17][20],S[149],C[149]);
  fa FA_00000150 (P[18][19],P[19][18],P[20][17],S[150],C[150]);
  fa FA_00000151 (P[21][16],P[22][15],P[23][14],S[151],C[151]);
  fa FA_00000152 (P[24][13],P[25][12],P[26][11],S[152],C[152]);
  fa FA_00000153 (P[27][10],P[28][9],P[29][8],S[153],C[153]);
  fa FA_00000154 (P[7][31],P[8][30],P[9][29],S[154],C[154]);
  fa FA_00000155 (P[10][28],P[11][27],P[12][26],S[155],C[155]);
  fa FA_00000156 (P[13][25],P[14][24],P[15][23],S[156],C[156]);
  fa FA_00000157 (P[16][22],P[17][21],P[18][20],S[157],C[157]);
  fa FA_00000158 (P[19][19],P[20][18],P[21][17],S[158],C[158]);
  fa FA_00000159 (P[22][16],P[23][15],P[24][14],S[159],C[159]);
  fa FA_00000160 (P[25][13],P[26][12],P[27][11],S[160],C[160]);
  fa FA_00000161 (P[8][31],P[9][30],P[10][29],S[161],C[161]);
  fa FA_00000162 (P[11][28],P[12][27],P[13][26],S[162],C[162]);
  fa FA_00000163 (P[14][25],P[15][24],P[16][23],S[163],C[163]);
  fa FA_00000164 (P[17][22],P[18][21],P[19][20],S[164],C[164]);
  fa FA_00000165 (P[20][19],P[21][18],P[22][17],S[165],C[165]);
  fa FA_00000166 (P[23][16],P[24][15],P[25][14],S[166],C[166]);
  fa FA_00000167 (P[9][31],P[10][30],P[11][29],S[167],C[167]);
  fa FA_00000168 (P[12][28],P[13][27],P[14][26],S[168],C[168]);
  fa FA_00000169 (P[15][25],P[16][24],P[17][23],S[169],C[169]);
  fa FA_00000170 (P[18][22],P[19][21],P[20][20],S[170],C[170]);
  fa FA_00000171 (P[21][19],P[22][18],P[23][17],S[171],C[171]);
  fa FA_00000172 (P[10][31],P[11][30],P[12][29],S[172],C[172]);
  fa FA_00000173 (P[13][28],P[14][27],P[15][26],S[173],C[173]);
  fa FA_00000174 (P[16][25],P[17][24],P[18][23],S[174],C[174]);
  fa FA_00000175 (P[19][22],P[20][21],P[21][20],S[175],C[175]);
  fa FA_00000176 (P[11][31],P[12][30],P[13][29],S[176],C[176]);
  fa FA_00000177 (P[14][28],P[15][27],P[16][26],S[177],C[177]);
  fa FA_00000178 (P[17][25],P[18][24],P[19][23],S[178],C[178]);
  fa FA_00000179 (P[12][31],P[13][30],P[14][29],S[179],C[179]);
  fa FA_00000180 (P[15][28],P[16][27],P[17][26],S[180],C[180]);
  fa FA_00000181 (P[13][31],P[14][30],P[15][29],S[181],C[181]);
  ha HA_00000182 (P[0][13],P[1][12],S[182],C[182]);
  fa FA_00000183 (P[0][14],P[1][13],P[2][12],S[183],C[183]);
  ha HA_00000184 (P[3][11],P[4][10],S[184],C[184]);
  fa FA_00000185 (P[0][15],P[1][14],P[2][13],S[185],C[185]);
  fa FA_00000186 (P[3][12],P[4][11],P[5][10],S[186],C[186]);
  ha HA_00000187 (P[6][9],P[7][8],S[187],C[187]);
  fa FA_00000188 (P[0][16],P[1][15],P[2][14],S[188],C[188]);
  fa FA_00000189 (P[3][13],P[4][12],P[5][11],S[189],C[189]);
  fa FA_00000190 (P[6][10],P[7][9],P[8][8],S[190],C[190]);
  ha HA_00000191 (P[9][7],P[10][6],S[191],C[191]);
  fa FA_00000192 (P[0][17],P[1][16],P[2][15],S[192],C[192]);
  fa FA_00000193 (P[3][14],P[4][13],P[5][12],S[193],C[193]);
  fa FA_00000194 (P[6][11],P[7][10],P[8][9],S[194],C[194]);
  fa FA_00000195 (P[9][8],P[10][7],P[11][6],S[195],C[195]);
  ha HA_00000196 (P[12][5],P[13][4],S[196],C[196]);
  fa FA_00000197 (P[0][18],P[1][17],P[2][16],S[197],C[197]);
  fa FA_00000198 (P[3][15],P[4][14],P[5][13],S[198],C[198]);
  fa FA_00000199 (P[6][12],P[7][11],P[8][10],S[199],C[199]);
  fa FA_00000200 (P[9][9],P[10][8],P[11][7],S[200],C[200]);
  fa FA_00000201 (P[12][6],P[13][5],P[14][4],S[201],C[201]);
  ha HA_00000202 (P[15][3],P[16][2],S[202],C[202]);
  fa FA_00000203 (S[20],P[2][17],P[3][16],S[203],C[203]);
  fa FA_00000204 (P[4][15],P[5][14],P[6][13],S[204],C[204]);
  fa FA_00000205 (P[7][12],P[8][11],P[9][10],S[205],C[205]);
  fa FA_00000206 (P[10][9],P[11][8],P[12][7],S[206],C[206]);
  fa FA_00000207 (P[13][6],P[14][5],P[15][4],S[207],C[207]);
  fa FA_00000208 (P[16][3],P[17][2],P[18][1],S[208],C[208]);
  fa FA_00000209 (S[21],C[20],S[22],S[209],C[209]);
  fa FA_00000210 (P[5][15],P[6][14],P[7][13],S[210],C[210]);
  fa FA_00000211 (P[8][12],P[9][11],P[10][10],S[211],C[211]);
  fa FA_00000212 (P[11][9],P[12][8],P[13][7],S[212],C[212]);
  fa FA_00000213 (P[14][6],P[15][5],P[16][4],S[213],C[213]);
  fa FA_00000214 (P[17][3],P[18][2],P[19][1],S[214],C[214]);
  fa FA_00000215 (S[23],C[21],S[24],S[215],C[215]);
  fa FA_00000216 (C[22],S[25],P[8][13],S[216],C[216]);
  fa FA_00000217 (P[9][12],P[10][11],P[11][10],S[217],C[217]);
  fa FA_00000218 (P[12][9],P[13][8],P[14][7],S[218],C[218]);
  fa FA_00000219 (P[15][6],P[16][5],P[17][4],S[219],C[219]);
  fa FA_00000220 (P[18][3],P[19][2],P[20][1],S[220],C[220]);
  fa FA_00000221 (S[26],C[23],S[27],S[221],C[221]);
  fa FA_00000222 (C[24],S[28],C[25],S[222],C[222]);
  fa FA_00000223 (S[29],P[11][11],P[12][10],S[223],C[223]);
  fa FA_00000224 (P[13][9],P[14][8],P[15][7],S[224],C[224]);
  fa FA_00000225 (P[16][6],P[17][5],P[18][4],S[225],C[225]);
  fa FA_00000226 (P[19][3],P[20][2],P[21][1],S[226],C[226]);
  fa FA_00000227 (S[30],C[26],S[31],S[227],C[227]);
  fa FA_00000228 (C[27],S[32],C[28],S[228],C[228]);
  fa FA_00000229 (S[33],C[29],S[34],S[229],C[229]);
  fa FA_00000230 (P[14][9],P[15][8],P[16][7],S[230],C[230]);
  fa FA_00000231 (P[17][6],P[18][5],P[19][4],S[231],C[231]);
  fa FA_00000232 (P[20][3],P[21][2],P[22][1],S[232],C[232]);
  fa FA_00000233 (S[35],C[30],S[36],S[233],C[233]);
  fa FA_00000234 (C[31],S[37],C[32],S[234],C[234]);
  fa FA_00000235 (S[38],C[33],S[39],S[235],C[235]);
  fa FA_00000236 (C[34],S[40],P[17][7],S[236],C[236]);
  fa FA_00000237 (P[18][6],P[19][5],P[20][4],S[237],C[237]);
  fa FA_00000238 (P[21][3],P[22][2],P[23][1],S[238],C[238]);
  fa FA_00000239 (S[41],C[35],S[42],S[239],C[239]);
  fa FA_00000240 (C[36],S[43],C[37],S[240],C[240]);
  fa FA_00000241 (S[44],C[38],S[45],S[241],C[241]);
  fa FA_00000242 (C[39],S[46],C[40],S[242],C[242]);
  fa FA_00000243 (S[47],P[20][5],P[21][4],S[243],C[243]);
  fa FA_00000244 (P[22][3],P[23][2],P[24][1],S[244],C[244]);
  fa FA_00000245 (S[48],C[41],S[49],S[245],C[245]);
  fa FA_00000246 (C[42],S[50],C[43],S[246],C[246]);
  fa FA_00000247 (S[51],C[44],S[52],S[247],C[247]);
  fa FA_00000248 (C[45],S[53],C[46],S[248],C[248]);
  fa FA_00000249 (S[54],C[47],S[55],S[249],C[249]);
  fa FA_00000250 (P[23][3],P[24][2],P[25][1],S[250],C[250]);
  fa FA_00000251 (S[56],C[48],S[57],S[251],C[251]);
  fa FA_00000252 (C[49],S[58],C[50],S[252],C[252]);
  fa FA_00000253 (S[59],C[51],S[60],S[253],C[253]);
  fa FA_00000254 (C[52],S[61],C[53],S[254],C[254]);
  fa FA_00000255 (S[62],C[54],S[63],S[255],C[255]);
  fa FA_00000256 (C[55],S[64],P[26][1],S[256],C[256]);
  fa FA_00000257 (S[65],C[56],S[66],S[257],C[257]);
  fa FA_00000258 (C[57],S[67],C[58],S[258],C[258]);
  fa FA_00000259 (S[68],C[59],S[69],S[259],C[259]);
  fa FA_00000260 (C[60],S[70],C[61],S[260],C[260]);
  fa FA_00000261 (S[71],C[62],S[72],S[261],C[261]);
  fa FA_00000262 (C[63],S[73],C[64],S[262],C[262]);
  fa FA_00000263 (S[74],C[65],S[75],S[263],C[263]);
  fa FA_00000264 (C[66],S[76],C[67],S[264],C[264]);
  fa FA_00000265 (S[77],C[68],S[78],S[265],C[265]);
  fa FA_00000266 (C[69],S[79],C[70],S[266],C[266]);
  fa FA_00000267 (S[80],C[71],S[81],S[267],C[267]);
  fa FA_00000268 (C[72],S[82],C[73],S[268],C[268]);
  fa FA_00000269 (S[83],C[74],S[84],S[269],C[269]);
  fa FA_00000270 (C[75],S[85],C[76],S[270],C[270]);
  fa FA_00000271 (S[86],C[77],S[87],S[271],C[271]);
  fa FA_00000272 (C[78],S[88],C[79],S[272],C[272]);
  fa FA_00000273 (S[89],C[80],S[90],S[273],C[273]);
  fa FA_00000274 (C[81],S[91],C[82],S[274],C[274]);
  fa FA_00000275 (S[92],C[83],S[93],S[275],C[275]);
  fa FA_00000276 (C[84],S[94],C[85],S[276],C[276]);
  fa FA_00000277 (S[95],C[86],S[96],S[277],C[277]);
  fa FA_00000278 (C[87],S[97],C[88],S[278],C[278]);
  fa FA_00000279 (S[98],C[89],S[99],S[279],C[279]);
  fa FA_00000280 (C[90],S[100],C[91],S[280],C[280]);
  fa FA_00000281 (S[101],C[92],S[102],S[281],C[281]);
  fa FA_00000282 (C[93],S[103],C[94],S[282],C[282]);
  fa FA_00000283 (S[104],C[95],S[105],S[283],C[283]);
  fa FA_00000284 (C[96],S[106],C[97],S[284],C[284]);
  fa FA_00000285 (S[107],C[98],S[108],S[285],C[285]);
  fa FA_00000286 (C[99],S[109],C[100],S[286],C[286]);
  fa FA_00000287 (S[110],C[101],S[111],S[287],C[287]);
  fa FA_00000288 (C[102],S[112],C[103],S[288],C[288]);
  fa FA_00000289 (S[113],C[104],S[114],S[289],C[289]);
  fa FA_00000290 (C[105],S[115],C[106],S[290],C[290]);
  fa FA_00000291 (S[116],C[107],S[117],S[291],C[291]);
  fa FA_00000292 (C[108],S[118],C[109],S[292],C[292]);
  fa FA_00000293 (S[119],C[110],S[120],S[293],C[293]);
  fa FA_00000294 (C[111],S[121],C[112],S[294],C[294]);
  fa FA_00000295 (S[122],C[113],S[123],S[295],C[295]);
  fa FA_00000296 (C[114],S[124],C[115],S[296],C[296]);
  fa FA_00000297 (S[125],C[116],S[126],S[297],C[297]);
  fa FA_00000298 (C[117],S[127],C[118],S[298],C[298]);
  fa FA_00000299 (S[128],C[119],S[129],S[299],C[299]);
  fa FA_00000300 (C[120],S[130],C[121],S[300],C[300]);
  fa FA_00000301 (S[131],C[122],S[132],S[301],C[301]);
  fa FA_00000302 (C[123],S[133],C[124],S[302],C[302]);
  fa FA_00000303 (S[134],C[125],S[135],S[303],C[303]);
  fa FA_00000304 (C[126],S[136],C[127],S[304],C[304]);
  fa FA_00000305 (S[137],C[128],S[138],S[305],C[305]);
  fa FA_00000306 (C[129],S[139],C[130],S[306],C[306]);
  fa FA_00000307 (S[140],C[131],S[141],S[307],C[307]);
  fa FA_00000308 (C[132],S[142],C[133],S[308],C[308]);
  fa FA_00000309 (S[143],C[134],S[144],S[309],C[309]);
  fa FA_00000310 (C[135],S[145],C[136],S[310],C[310]);
  fa FA_00000311 (S[146],C[137],S[147],S[311],C[311]);
  fa FA_00000312 (C[138],S[148],C[139],S[312],C[312]);
  fa FA_00000313 (S[149],C[140],S[150],S[313],C[313]);
  fa FA_00000314 (C[141],S[151],C[142],S[314],C[314]);
  fa FA_00000315 (S[152],C[143],S[153],S[315],C[315]);
  fa FA_00000316 (C[144],C[145],P[30][7],S[316],C[316]);
  fa FA_00000317 (S[154],C[146],S[155],S[317],C[317]);
  fa FA_00000318 (C[147],S[156],C[148],S[318],C[318]);
  fa FA_00000319 (S[157],C[149],S[158],S[319],C[319]);
  fa FA_00000320 (C[150],S[159],C[151],S[320],C[320]);
  fa FA_00000321 (S[160],C[152],C[153],S[321],C[321]);
  fa FA_00000322 (P[28][10],P[29][9],P[30][8],S[322],C[322]);
  fa FA_00000323 (S[161],C[154],S[162],S[323],C[323]);
  fa FA_00000324 (C[155],S[163],C[156],S[324],C[324]);
  fa FA_00000325 (S[164],C[157],S[165],S[325],C[325]);
  fa FA_00000326 (C[158],S[166],C[159],S[326],C[326]);
  fa FA_00000327 (C[160],P[26][13],P[27][12],S[327],C[327]);
  fa FA_00000328 (P[28][11],P[29][10],P[30][9],S[328],C[328]);
  fa FA_00000329 (S[167],C[161],S[168],S[329],C[329]);
  fa FA_00000330 (C[162],S[169],C[163],S[330],C[330]);
  fa FA_00000331 (S[170],C[164],S[171],S[331],C[331]);
  fa FA_00000332 (C[165],C[166],P[24][16],S[332],C[332]);
  fa FA_00000333 (P[25][15],P[26][14],P[27][13],S[333],C[333]);
  fa FA_00000334 (P[28][12],P[29][11],P[30][10],S[334],C[334]);
  fa FA_00000335 (S[172],C[167],S[173],S[335],C[335]);
  fa FA_00000336 (C[168],S[174],C[169],S[336],C[336]);
  fa FA_00000337 (S[175],C[170],C[171],S[337],C[337]);
  fa FA_00000338 (P[22][19],P[23][18],P[24][17],S[338],C[338]);
  fa FA_00000339 (P[25][16],P[26][15],P[27][14],S[339],C[339]);
  fa FA_00000340 (P[28][13],P[29][12],P[30][11],S[340],C[340]);
  fa FA_00000341 (S[176],C[172],S[177],S[341],C[341]);
  fa FA_00000342 (C[173],S[178],C[174],S[342],C[342]);
  fa FA_00000343 (C[175],P[20][22],P[21][21],S[343],C[343]);
  fa FA_00000344 (P[22][20],P[23][19],P[24][18],S[344],C[344]);
  fa FA_00000345 (P[25][17],P[26][16],P[27][15],S[345],C[345]);
  fa FA_00000346 (P[28][14],P[29][13],P[30][12],S[346],C[346]);
  fa FA_00000347 (S[179],C[176],S[180],S[347],C[347]);
  fa FA_00000348 (C[177],C[178],P[18][25],S[348],C[348]);
  fa FA_00000349 (P[19][24],P[20][23],P[21][22],S[349],C[349]);
  fa FA_00000350 (P[22][21],P[23][20],P[24][19],S[350],C[350]);
  fa FA_00000351 (P[25][18],P[26][17],P[27][16],S[351],C[351]);
  fa FA_00000352 (P[28][15],P[29][14],P[30][13],S[352],C[352]);
  fa FA_00000353 (S[181],C[179],C[180],S[353],C[353]);
  fa FA_00000354 (P[16][28],P[17][27],P[18][26],S[354],C[354]);
  fa FA_00000355 (P[19][25],P[20][24],P[21][23],S[355],C[355]);
  fa FA_00000356 (P[22][22],P[23][21],P[24][20],S[356],C[356]);
  fa FA_00000357 (P[25][19],P[26][18],P[27][17],S[357],C[357]);
  fa FA_00000358 (P[28][16],P[29][15],P[30][14],S[358],C[358]);
  fa FA_00000359 (C[181],P[14][31],P[15][30],S[359],C[359]);
  fa FA_00000360 (P[16][29],P[17][28],P[18][27],S[360],C[360]);
  fa FA_00000361 (P[19][26],P[20][25],P[21][24],S[361],C[361]);
  fa FA_00000362 (P[22][23],P[23][22],P[24][21],S[362],C[362]);
  fa FA_00000363 (P[25][20],P[26][19],P[27][18],S[363],C[363]);
  fa FA_00000364 (P[28][17],P[29][16],P[30][15],S[364],C[364]);
  fa FA_00000365 (P[15][31],P[16][30],P[17][29],S[365],C[365]);
  fa FA_00000366 (P[18][28],P[19][27],P[20][26],S[366],C[366]);
  fa FA_00000367 (P[21][25],P[22][24],P[23][23],S[367],C[367]);
  fa FA_00000368 (P[24][22],P[25][21],P[26][20],S[368],C[368]);
  fa FA_00000369 (P[27][19],P[28][18],P[29][17],S[369],C[369]);
  fa FA_00000370 (P[16][31],P[17][30],P[18][29],S[370],C[370]);
  fa FA_00000371 (P[19][28],P[20][27],P[21][26],S[371],C[371]);
  fa FA_00000372 (P[22][25],P[23][24],P[24][23],S[372],C[372]);
  fa FA_00000373 (P[25][22],P[26][21],P[27][20],S[373],C[373]);
  fa FA_00000374 (P[17][31],P[18][30],P[19][29],S[374],C[374]);
  fa FA_00000375 (P[20][28],P[21][27],P[22][26],S[375],C[375]);
  fa FA_00000376 (P[23][25],P[24][24],P[25][23],S[376],C[376]);
  fa FA_00000377 (P[18][31],P[19][30],P[20][29],S[377],C[377]);
  fa FA_00000378 (P[21][28],P[22][27],P[23][26],S[378],C[378]);
  fa FA_00000379 (P[19][31],P[20][30],P[21][29],S[379],C[379]);
  ha HA_00000380 (P[0][9],P[1][8],S[380],C[380]);
  fa FA_00000381 (P[0][10],P[1][9],P[2][8],S[381],C[381]);
  ha HA_00000382 (P[3][7],P[4][6],S[382],C[382]);
  fa FA_00000383 (P[0][11],P[1][10],P[2][9],S[383],C[383]);
  fa FA_00000384 (P[3][8],P[4][7],P[5][6],S[384],C[384]);
  ha HA_00000385 (P[6][5],P[7][4],S[385],C[385]);
  fa FA_00000386 (P[0][12],P[1][11],P[2][10],S[386],C[386]);
  fa FA_00000387 (P[3][9],P[4][8],P[5][7],S[387],C[387]);
  fa FA_00000388 (P[6][6],P[7][5],P[8][4],S[388],C[388]);
  ha HA_00000389 (P[9][3],P[10][2],S[389],C[389]);
  fa FA_00000390 (S[182],P[2][11],P[3][10],S[390],C[390]);
  fa FA_00000391 (P[4][9],P[5][8],P[6][7],S[391],C[391]);
  fa FA_00000392 (P[7][6],P[8][5],P[9][4],S[392],C[392]);
  fa FA_00000393 (P[10][3],P[11][2],P[12][1],S[393],C[393]);
  fa FA_00000394 (S[183],C[182],S[184],S[394],C[394]);
  fa FA_00000395 (P[5][9],P[6][8],P[7][7],S[395],C[395]);
  fa FA_00000396 (P[8][6],P[9][5],P[10][4],S[396],C[396]);
  fa FA_00000397 (P[11][3],P[12][2],P[13][1],S[397],C[397]);
  fa FA_00000398 (S[185],C[183],S[186],S[398],C[398]);
  fa FA_00000399 (C[184],S[187],P[8][7],S[399],C[399]);
  fa FA_00000400 (P[9][6],P[10][5],P[11][4],S[400],C[400]);
  fa FA_00000401 (P[12][3],P[13][2],P[14][1],S[401],C[401]);
  fa FA_00000402 (S[188],C[185],S[189],S[402],C[402]);
  fa FA_00000403 (C[186],S[190],C[187],S[403],C[403]);
  fa FA_00000404 (S[191],P[11][5],P[12][4],S[404],C[404]);
  fa FA_00000405 (P[13][3],P[14][2],P[15][1],S[405],C[405]);
  fa FA_00000406 (S[192],C[188],S[193],S[406],C[406]);
  fa FA_00000407 (C[189],S[194],C[190],S[407],C[407]);
  fa FA_00000408 (S[195],C[191],S[196],S[408],C[408]);
  fa FA_00000409 (P[14][3],P[15][2],P[16][1],S[409],C[409]);
  fa FA_00000410 (S[197],C[192],S[198],S[410],C[410]);
  fa FA_00000411 (C[193],S[199],C[194],S[411],C[411]);
  fa FA_00000412 (S[200],C[195],S[201],S[412],C[412]);
  fa FA_00000413 (C[196],S[202],P[17][1],S[413],C[413]);
  fa FA_00000414 (S[203],C[197],S[204],S[414],C[414]);
  fa FA_00000415 (C[198],S[205],C[199],S[415],C[415]);
  fa FA_00000416 (S[206],C[200],S[207],S[416],C[416]);
  fa FA_00000417 (C[201],S[208],C[202],S[417],C[417]);
  fa FA_00000418 (S[209],C[203],S[210],S[418],C[418]);
  fa FA_00000419 (C[204],S[211],C[205],S[419],C[419]);
  fa FA_00000420 (S[212],C[206],S[213],S[420],C[420]);
  fa FA_00000421 (C[207],S[214],C[208],S[421],C[421]);
  fa FA_00000422 (S[215],C[209],S[216],S[422],C[422]);
  fa FA_00000423 (C[210],S[217],C[211],S[423],C[423]);
  fa FA_00000424 (S[218],C[212],S[219],S[424],C[424]);
  fa FA_00000425 (C[213],S[220],C[214],S[425],C[425]);
  fa FA_00000426 (S[221],C[215],S[222],S[426],C[426]);
  fa FA_00000427 (C[216],S[223],C[217],S[427],C[427]);
  fa FA_00000428 (S[224],C[218],S[225],S[428],C[428]);
  fa FA_00000429 (C[219],S[226],C[220],S[429],C[429]);
  fa FA_00000430 (S[227],C[221],S[228],S[430],C[430]);
  fa FA_00000431 (C[222],S[229],C[223],S[431],C[431]);
  fa FA_00000432 (S[230],C[224],S[231],S[432],C[432]);
  fa FA_00000433 (C[225],S[232],C[226],S[433],C[433]);
  fa FA_00000434 (S[233],C[227],S[234],S[434],C[434]);
  fa FA_00000435 (C[228],S[235],C[229],S[435],C[435]);
  fa FA_00000436 (S[236],C[230],S[237],S[436],C[436]);
  fa FA_00000437 (C[231],S[238],C[232],S[437],C[437]);
  fa FA_00000438 (S[239],C[233],S[240],S[438],C[438]);
  fa FA_00000439 (C[234],S[241],C[235],S[439],C[439]);
  fa FA_00000440 (S[242],C[236],S[243],S[440],C[440]);
  fa FA_00000441 (C[237],S[244],C[238],S[441],C[441]);
  fa FA_00000442 (S[245],C[239],S[246],S[442],C[442]);
  fa FA_00000443 (C[240],S[247],C[241],S[443],C[443]);
  fa FA_00000444 (S[248],C[242],S[249],S[444],C[444]);
  fa FA_00000445 (C[243],S[250],C[244],S[445],C[445]);
  fa FA_00000446 (S[251],C[245],S[252],S[446],C[446]);
  fa FA_00000447 (C[246],S[253],C[247],S[447],C[447]);
  fa FA_00000448 (S[254],C[248],S[255],S[448],C[448]);
  fa FA_00000449 (C[249],S[256],C[250],S[449],C[449]);
  fa FA_00000450 (S[257],C[251],S[258],S[450],C[450]);
  fa FA_00000451 (C[252],S[259],C[253],S[451],C[451]);
  fa FA_00000452 (S[260],C[254],S[261],S[452],C[452]);
  fa FA_00000453 (C[255],S[262],C[256],S[453],C[453]);
  fa FA_00000454 (S[263],C[257],S[264],S[454],C[454]);
  fa FA_00000455 (C[258],S[265],C[259],S[455],C[455]);
  fa FA_00000456 (S[266],C[260],S[267],S[456],C[456]);
  fa FA_00000457 (C[261],S[268],C[262],S[457],C[457]);
  fa FA_00000458 (S[269],C[263],S[270],S[458],C[458]);
  fa FA_00000459 (C[264],S[271],C[265],S[459],C[459]);
  fa FA_00000460 (S[272],C[266],S[273],S[460],C[460]);
  fa FA_00000461 (C[267],S[274],C[268],S[461],C[461]);
  fa FA_00000462 (S[275],C[269],S[276],S[462],C[462]);
  fa FA_00000463 (C[270],S[277],C[271],S[463],C[463]);
  fa FA_00000464 (S[278],C[272],S[279],S[464],C[464]);
  fa FA_00000465 (C[273],S[280],C[274],S[465],C[465]);
  fa FA_00000466 (S[281],C[275],S[282],S[466],C[466]);
  fa FA_00000467 (C[276],S[283],C[277],S[467],C[467]);
  fa FA_00000468 (S[284],C[278],S[285],S[468],C[468]);
  fa FA_00000469 (C[279],S[286],C[280],S[469],C[469]);
  fa FA_00000470 (S[287],C[281],S[288],S[470],C[470]);
  fa FA_00000471 (C[282],S[289],C[283],S[471],C[471]);
  fa FA_00000472 (S[290],C[284],S[291],S[472],C[472]);
  fa FA_00000473 (C[285],S[292],C[286],S[473],C[473]);
  fa FA_00000474 (S[293],C[287],S[294],S[474],C[474]);
  fa FA_00000475 (C[288],S[295],C[289],S[475],C[475]);
  fa FA_00000476 (S[296],C[290],S[297],S[476],C[476]);
  fa FA_00000477 (C[291],S[298],C[292],S[477],C[477]);
  fa FA_00000478 (S[299],C[293],S[300],S[478],C[478]);
  fa FA_00000479 (C[294],S[301],C[295],S[479],C[479]);
  fa FA_00000480 (S[302],C[296],S[303],S[480],C[480]);
  fa FA_00000481 (C[297],S[304],C[298],S[481],C[481]);
  fa FA_00000482 (S[305],C[299],S[306],S[482],C[482]);
  fa FA_00000483 (C[300],S[307],C[301],S[483],C[483]);
  fa FA_00000484 (S[308],C[302],S[309],S[484],C[484]);
  fa FA_00000485 (C[303],S[310],C[304],S[485],C[485]);
  fa FA_00000486 (S[311],C[305],S[312],S[486],C[486]);
  fa FA_00000487 (C[306],S[313],C[307],S[487],C[487]);
  fa FA_00000488 (S[314],C[308],S[315],S[488],C[488]);
  fa FA_00000489 (C[309],S[316],C[310],S[489],C[489]);
  fa FA_00000490 (S[317],C[311],S[318],S[490],C[490]);
  fa FA_00000491 (C[312],S[319],C[313],S[491],C[491]);
  fa FA_00000492 (S[320],C[314],S[321],S[492],C[492]);
  fa FA_00000493 (C[315],S[322],C[316],S[493],C[493]);
  fa FA_00000494 (S[323],C[317],S[324],S[494],C[494]);
  fa FA_00000495 (C[318],S[325],C[319],S[495],C[495]);
  fa FA_00000496 (S[326],C[320],S[327],S[496],C[496]);
  fa FA_00000497 (C[321],S[328],C[322],S[497],C[497]);
  fa FA_00000498 (S[329],C[323],S[330],S[498],C[498]);
  fa FA_00000499 (C[324],S[331],C[325],S[499],C[499]);
  fa FA_00000500 (S[332],C[326],S[333],S[500],C[500]);
  fa FA_00000501 (C[327],S[334],C[328],S[501],C[501]);
  fa FA_00000502 (S[335],C[329],S[336],S[502],C[502]);
  fa FA_00000503 (C[330],S[337],C[331],S[503],C[503]);
  fa FA_00000504 (S[338],C[332],S[339],S[504],C[504]);
  fa FA_00000505 (C[333],S[340],C[334],S[505],C[505]);
  fa FA_00000506 (S[341],C[335],S[342],S[506],C[506]);
  fa FA_00000507 (C[336],S[343],C[337],S[507],C[507]);
  fa FA_00000508 (S[344],C[338],S[345],S[508],C[508]);
  fa FA_00000509 (C[339],S[346],C[340],S[509],C[509]);
  fa FA_00000510 (S[347],C[341],S[348],S[510],C[510]);
  fa FA_00000511 (C[342],S[349],C[343],S[511],C[511]);
  fa FA_00000512 (S[350],C[344],S[351],S[512],C[512]);
  fa FA_00000513 (C[345],S[352],C[346],S[513],C[513]);
  fa FA_00000514 (S[353],C[347],S[354],S[514],C[514]);
  fa FA_00000515 (C[348],S[355],C[349],S[515],C[515]);
  fa FA_00000516 (S[356],C[350],S[357],S[516],C[516]);
  fa FA_00000517 (C[351],S[358],C[352],S[517],C[517]);
  fa FA_00000518 (S[359],C[353],S[360],S[518],C[518]);
  fa FA_00000519 (C[354],S[361],C[355],S[519],C[519]);
  fa FA_00000520 (S[362],C[356],S[363],S[520],C[520]);
  fa FA_00000521 (C[357],S[364],C[358],S[521],C[521]);
  fa FA_00000522 (S[365],C[359],S[366],S[522],C[522]);
  fa FA_00000523 (C[360],S[367],C[361],S[523],C[523]);
  fa FA_00000524 (S[368],C[362],S[369],S[524],C[524]);
  fa FA_00000525 (C[363],C[364],P[30][16],S[525],C[525]);
  fa FA_00000526 (S[370],C[365],S[371],S[526],C[526]);
  fa FA_00000527 (C[366],S[372],C[367],S[527],C[527]);
  fa FA_00000528 (S[373],C[368],C[369],S[528],C[528]);
  fa FA_00000529 (P[28][19],P[29][18],P[30][17],S[529],C[529]);
  fa FA_00000530 (S[374],C[370],S[375],S[530],C[530]);
  fa FA_00000531 (C[371],S[376],C[372],S[531],C[531]);
  fa FA_00000532 (C[373],P[26][22],P[27][21],S[532],C[532]);
  fa FA_00000533 (P[28][20],P[29][19],P[30][18],S[533],C[533]);
  fa FA_00000534 (S[377],C[374],S[378],S[534],C[534]);
  fa FA_00000535 (C[375],C[376],P[24][25],S[535],C[535]);
  fa FA_00000536 (P[25][24],P[26][23],P[27][22],S[536],C[536]);
  fa FA_00000537 (P[28][21],P[29][20],P[30][19],S[537],C[537]);
  fa FA_00000538 (S[379],C[377],C[378],S[538],C[538]);
  fa FA_00000539 (P[22][28],P[23][27],P[24][26],S[539],C[539]);
  fa FA_00000540 (P[25][25],P[26][24],P[27][23],S[540],C[540]);
  fa FA_00000541 (P[28][22],P[29][21],P[30][20],S[541],C[541]);
  fa FA_00000542 (C[379],P[20][31],P[21][30],S[542],C[542]);
  fa FA_00000543 (P[22][29],P[23][28],P[24][27],S[543],C[543]);
  fa FA_00000544 (P[25][26],P[26][25],P[27][24],S[544],C[544]);
  fa FA_00000545 (P[28][23],P[29][22],P[30][21],S[545],C[545]);
  fa FA_00000546 (P[21][31],P[22][30],P[23][29],S[546],C[546]);
  fa FA_00000547 (P[24][28],P[25][27],P[26][26],S[547],C[547]);
  fa FA_00000548 (P[27][25],P[28][24],P[29][23],S[548],C[548]);
  fa FA_00000549 (P[22][31],P[23][30],P[24][29],S[549],C[549]);
  fa FA_00000550 (P[25][28],P[26][27],P[27][26],S[550],C[550]);
  fa FA_00000551 (P[23][31],P[24][30],P[25][29],S[551],C[551]);
  ha HA_00000552 (P[0][6],P[1][5],S[552],C[552]);
  fa FA_00000553 (P[0][7],P[1][6],P[2][5],S[553],C[553]);
  ha HA_00000554 (P[3][4],P[4][3],S[554],C[554]);
  fa FA_00000555 (P[0][8],P[1][7],P[2][6],S[555],C[555]);
  fa FA_00000556 (P[3][5],P[4][4],P[5][3],S[556],C[556]);
  ha HA_00000557 (P[6][2],P[7][1],S[557],C[557]);
  fa FA_00000558 (S[380],P[2][7],P[3][6],S[558],C[558]);
  fa FA_00000559 (P[4][5],P[5][4],P[6][3],S[559],C[559]);
  fa FA_00000560 (P[7][2],P[8][1],P[9][0],S[560],C[560]);
  fa FA_00000561 (S[381],C[380],S[382],S[561],C[561]);
  fa FA_00000562 (P[5][5],P[6][4],P[7][3],S[562],C[562]);
  fa FA_00000563 (P[8][2],P[9][1],P[10][0],S[563],C[563]);
  fa FA_00000564 (S[383],C[381],S[384],S[564],C[564]);
  fa FA_00000565 (C[382],S[385],P[8][3],S[565],C[565]);
  fa FA_00000566 (P[9][2],P[10][1],P[11][0],S[566],C[566]);
  fa FA_00000567 (S[386],C[383],S[387],S[567],C[567]);
  fa FA_00000568 (C[384],S[388],C[385],S[568],C[568]);
  fa FA_00000569 (S[389],P[11][1],P[12][0],S[569],C[569]);
  fa FA_00000570 (S[390],C[386],S[391],S[570],C[570]);
  fa FA_00000571 (C[387],S[392],C[388],S[571],C[571]);
  fa FA_00000572 (S[393],C[389],P[13][0],S[572],C[572]);
  fa FA_00000573 (S[394],C[390],S[395],S[573],C[573]);
  fa FA_00000574 (C[391],S[396],C[392],S[574],C[574]);
  fa FA_00000575 (S[397],C[393],P[14][0],S[575],C[575]);
  fa FA_00000576 (S[398],C[394],S[399],S[576],C[576]);
  fa FA_00000577 (C[395],S[400],C[396],S[577],C[577]);
  fa FA_00000578 (S[401],C[397],P[15][0],S[578],C[578]);
  fa FA_00000579 (S[402],C[398],S[403],S[579],C[579]);
  fa FA_00000580 (C[399],S[404],C[400],S[580],C[580]);
  fa FA_00000581 (S[405],C[401],P[16][0],S[581],C[581]);
  fa FA_00000582 (S[406],C[402],S[407],S[582],C[582]);
  fa FA_00000583 (C[403],S[408],C[404],S[583],C[583]);
  fa FA_00000584 (S[409],C[405],P[17][0],S[584],C[584]);
  fa FA_00000585 (S[410],C[406],S[411],S[585],C[585]);
  fa FA_00000586 (C[407],S[412],C[408],S[586],C[586]);
  fa FA_00000587 (S[413],C[409],P[18][0],S[587],C[587]);
  fa FA_00000588 (S[414],C[410],S[415],S[588],C[588]);
  fa FA_00000589 (C[411],S[416],C[412],S[589],C[589]);
  fa FA_00000590 (S[417],C[413],P[19][0],S[590],C[590]);
  fa FA_00000591 (S[418],C[414],S[419],S[591],C[591]);
  fa FA_00000592 (C[415],S[420],C[416],S[592],C[592]);
  fa FA_00000593 (S[421],C[417],P[20][0],S[593],C[593]);
  fa FA_00000594 (S[422],C[418],S[423],S[594],C[594]);
  fa FA_00000595 (C[419],S[424],C[420],S[595],C[595]);
  fa FA_00000596 (S[425],C[421],P[21][0],S[596],C[596]);
  fa FA_00000597 (S[426],C[422],S[427],S[597],C[597]);
  fa FA_00000598 (C[423],S[428],C[424],S[598],C[598]);
  fa FA_00000599 (S[429],C[425],P[22][0],S[599],C[599]);
  fa FA_00000600 (S[430],C[426],S[431],S[600],C[600]);
  fa FA_00000601 (C[427],S[432],C[428],S[601],C[601]);
  fa FA_00000602 (S[433],C[429],P[23][0],S[602],C[602]);
  fa FA_00000603 (S[434],C[430],S[435],S[603],C[603]);
  fa FA_00000604 (C[431],S[436],C[432],S[604],C[604]);
  fa FA_00000605 (S[437],C[433],P[24][0],S[605],C[605]);
  fa FA_00000606 (S[438],C[434],S[439],S[606],C[606]);
  fa FA_00000607 (C[435],S[440],C[436],S[607],C[607]);
  fa FA_00000608 (S[441],C[437],P[25][0],S[608],C[608]);
  fa FA_00000609 (S[442],C[438],S[443],S[609],C[609]);
  fa FA_00000610 (C[439],S[444],C[440],S[610],C[610]);
  fa FA_00000611 (S[445],C[441],P[26][0],S[611],C[611]);
  fa FA_00000612 (S[446],C[442],S[447],S[612],C[612]);
  fa FA_00000613 (C[443],S[448],C[444],S[613],C[613]);
  fa FA_00000614 (S[449],C[445],P[27][0],S[614],C[614]);
  fa FA_00000615 (S[450],C[446],S[451],S[615],C[615]);
  fa FA_00000616 (C[447],S[452],C[448],S[616],C[616]);
  fa FA_00000617 (S[453],C[449],P[28][0],S[617],C[617]);
  fa FA_00000618 (S[454],C[450],S[455],S[618],C[618]);
  fa FA_00000619 (C[451],S[456],C[452],S[619],C[619]);
  fa FA_00000620 (S[457],C[453],P[29][0],S[620],C[620]);
  fa FA_00000621 (S[458],C[454],S[459],S[621],C[621]);
  fa FA_00000622 (C[455],S[460],C[456],S[622],C[622]);
  fa FA_00000623 (S[461],C[457],P[30][0],S[623],C[623]);
  fa FA_00000624 (S[462],C[458],S[463],S[624],C[624]);
  fa FA_00000625 (C[459],S[464],C[460],S[625],C[625]);
  fa FA_00000626 (S[465],C[461],P[31][0],S[626],C[626]);
  fa FA_00000627 (S[466],C[462],S[467],S[627],C[627]);
  fa FA_00000628 (C[463],S[468],C[464],S[628],C[628]);
  fa FA_00000629 (S[469],C[465],P[31][1],S[629],C[629]);
  fa FA_00000630 (S[470],C[466],S[471],S[630],C[630]);
  fa FA_00000631 (C[467],S[472],C[468],S[631],C[631]);
  fa FA_00000632 (S[473],C[469],P[31][2],S[632],C[632]);
  fa FA_00000633 (S[474],C[470],S[475],S[633],C[633]);
  fa FA_00000634 (C[471],S[476],C[472],S[634],C[634]);
  fa FA_00000635 (S[477],C[473],P[31][3],S[635],C[635]);
  fa FA_00000636 (S[478],C[474],S[479],S[636],C[636]);
  fa FA_00000637 (C[475],S[480],C[476],S[637],C[637]);
  fa FA_00000638 (S[481],C[477],P[31][4],S[638],C[638]);
  fa FA_00000639 (S[482],C[478],S[483],S[639],C[639]);
  fa FA_00000640 (C[479],S[484],C[480],S[640],C[640]);
  fa FA_00000641 (S[485],C[481],P[31][5],S[641],C[641]);
  fa FA_00000642 (S[486],C[482],S[487],S[642],C[642]);
  fa FA_00000643 (C[483],S[488],C[484],S[643],C[643]);
  fa FA_00000644 (S[489],C[485],P[31][6],S[644],C[644]);
  fa FA_00000645 (S[490],C[486],S[491],S[645],C[645]);
  fa FA_00000646 (C[487],S[492],C[488],S[646],C[646]);
  fa FA_00000647 (S[493],C[489],P[31][7],S[647],C[647]);
  fa FA_00000648 (S[494],C[490],S[495],S[648],C[648]);
  fa FA_00000649 (C[491],S[496],C[492],S[649],C[649]);
  fa FA_00000650 (S[497],C[493],P[31][8],S[650],C[650]);
  fa FA_00000651 (S[498],C[494],S[499],S[651],C[651]);
  fa FA_00000652 (C[495],S[500],C[496],S[652],C[652]);
  fa FA_00000653 (S[501],C[497],P[31][9],S[653],C[653]);
  fa FA_00000654 (S[502],C[498],S[503],S[654],C[654]);
  fa FA_00000655 (C[499],S[504],C[500],S[655],C[655]);
  fa FA_00000656 (S[505],C[501],P[31][10],S[656],C[656]);
  fa FA_00000657 (S[506],C[502],S[507],S[657],C[657]);
  fa FA_00000658 (C[503],S[508],C[504],S[658],C[658]);
  fa FA_00000659 (S[509],C[505],P[31][11],S[659],C[659]);
  fa FA_00000660 (S[510],C[506],S[511],S[660],C[660]);
  fa FA_00000661 (C[507],S[512],C[508],S[661],C[661]);
  fa FA_00000662 (S[513],C[509],P[31][12],S[662],C[662]);
  fa FA_00000663 (S[514],C[510],S[515],S[663],C[663]);
  fa FA_00000664 (C[511],S[516],C[512],S[664],C[664]);
  fa FA_00000665 (S[517],C[513],P[31][13],S[665],C[665]);
  fa FA_00000666 (S[518],C[514],S[519],S[666],C[666]);
  fa FA_00000667 (C[515],S[520],C[516],S[667],C[667]);
  fa FA_00000668 (S[521],C[517],P[31][14],S[668],C[668]);
  fa FA_00000669 (S[522],C[518],S[523],S[669],C[669]);
  fa FA_00000670 (C[519],S[524],C[520],S[670],C[670]);
  fa FA_00000671 (S[525],C[521],P[31][15],S[671],C[671]);
  fa FA_00000672 (S[526],C[522],S[527],S[672],C[672]);
  fa FA_00000673 (C[523],S[528],C[524],S[673],C[673]);
  fa FA_00000674 (S[529],C[525],P[31][16],S[674],C[674]);
  fa FA_00000675 (S[530],C[526],S[531],S[675],C[675]);
  fa FA_00000676 (C[527],S[532],C[528],S[676],C[676]);
  fa FA_00000677 (S[533],C[529],P[31][17],S[677],C[677]);
  fa FA_00000678 (S[534],C[530],S[535],S[678],C[678]);
  fa FA_00000679 (C[531],S[536],C[532],S[679],C[679]);
  fa FA_00000680 (S[537],C[533],P[31][18],S[680],C[680]);
  fa FA_00000681 (S[538],C[534],S[539],S[681],C[681]);
  fa FA_00000682 (C[535],S[540],C[536],S[682],C[682]);
  fa FA_00000683 (S[541],C[537],P[31][19],S[683],C[683]);
  fa FA_00000684 (S[542],C[538],S[543],S[684],C[684]);
  fa FA_00000685 (C[539],S[544],C[540],S[685],C[685]);
  fa FA_00000686 (S[545],C[541],P[31][20],S[686],C[686]);
  fa FA_00000687 (S[546],C[542],S[547],S[687],C[687]);
  fa FA_00000688 (C[543],S[548],C[544],S[688],C[688]);
  fa FA_00000689 (C[545],P[30][22],P[31][21],S[689],C[689]);
  fa FA_00000690 (S[549],C[546],S[550],S[690],C[690]);
  fa FA_00000691 (C[547],C[548],P[28][25],S[691],C[691]);
  fa FA_00000692 (P[29][24],P[30][23],P[31][22],S[692],C[692]);
  fa FA_00000693 (S[551],C[549],C[550],S[693],C[693]);
  fa FA_00000694 (P[26][28],P[27][27],P[28][26],S[694],C[694]);
  fa FA_00000695 (P[29][25],P[30][24],P[31][23],S[695],C[695]);
  fa FA_00000696 (C[551],P[24][31],P[25][30],S[696],C[696]);
  fa FA_00000697 (P[26][29],P[27][28],P[28][27],S[697],C[697]);
  fa FA_00000698 (P[29][26],P[30][25],P[31][24],S[698],C[698]);
  fa FA_00000699 (P[25][31],P[26][30],P[27][29],S[699],C[699]);
  fa FA_00000700 (P[28][28],P[29][27],P[30][26],S[700],C[700]);
  fa FA_00000701 (P[26][31],P[27][30],P[28][29],S[701],C[701]);
  ha HA_00000702 (P[0][4],P[1][3],S[702],C[702]);
  fa FA_00000703 (P[0][5],P[1][4],P[2][3],S[703],C[703]);
  ha HA_00000704 (P[3][2],P[4][1],S[704],C[704]);
  fa FA_00000705 (S[552],P[2][4],P[3][3],S[705],C[705]);
  fa FA_00000706 (P[4][2],P[5][1],P[6][0],S[706],C[706]);
  fa FA_00000707 (S[553],C[552],S[554],S[707],C[707]);
  fa FA_00000708 (P[5][2],P[6][1],P[7][0],S[708],C[708]);
  fa FA_00000709 (S[555],C[553],S[556],S[709],C[709]);
  fa FA_00000710 (C[554],S[557],P[8][0],S[710],C[710]);
  fa FA_00000711 (S[558],C[555],S[559],S[711],C[711]);
  fa FA_00000712 (C[556],S[560],C[557],S[712],C[712]);
  fa FA_00000713 (S[561],C[558],S[562],S[713],C[713]);
  fa FA_00000714 (C[559],S[563],C[560],S[714],C[714]);
  fa FA_00000715 (S[564],C[561],S[565],S[715],C[715]);
  fa FA_00000716 (C[562],S[566],C[563],S[716],C[716]);
  fa FA_00000717 (S[567],C[564],S[568],S[717],C[717]);
  fa FA_00000718 (C[565],S[569],C[566],S[718],C[718]);
  fa FA_00000719 (S[570],C[567],S[571],S[719],C[719]);
  fa FA_00000720 (C[568],S[572],C[569],S[720],C[720]);
  fa FA_00000721 (S[573],C[570],S[574],S[721],C[721]);
  fa FA_00000722 (C[571],S[575],C[572],S[722],C[722]);
  fa FA_00000723 (S[576],C[573],S[577],S[723],C[723]);
  fa FA_00000724 (C[574],S[578],C[575],S[724],C[724]);
  fa FA_00000725 (S[579],C[576],S[580],S[725],C[725]);
  fa FA_00000726 (C[577],S[581],C[578],S[726],C[726]);
  fa FA_00000727 (S[582],C[579],S[583],S[727],C[727]);
  fa FA_00000728 (C[580],S[584],C[581],S[728],C[728]);
  fa FA_00000729 (S[585],C[582],S[586],S[729],C[729]);
  fa FA_00000730 (C[583],S[587],C[584],S[730],C[730]);
  fa FA_00000731 (S[588],C[585],S[589],S[731],C[731]);
  fa FA_00000732 (C[586],S[590],C[587],S[732],C[732]);
  fa FA_00000733 (S[591],C[588],S[592],S[733],C[733]);
  fa FA_00000734 (C[589],S[593],C[590],S[734],C[734]);
  fa FA_00000735 (S[594],C[591],S[595],S[735],C[735]);
  fa FA_00000736 (C[592],S[596],C[593],S[736],C[736]);
  fa FA_00000737 (S[597],C[594],S[598],S[737],C[737]);
  fa FA_00000738 (C[595],S[599],C[596],S[738],C[738]);
  fa FA_00000739 (S[600],C[597],S[601],S[739],C[739]);
  fa FA_00000740 (C[598],S[602],C[599],S[740],C[740]);
  fa FA_00000741 (S[603],C[600],S[604],S[741],C[741]);
  fa FA_00000742 (C[601],S[605],C[602],S[742],C[742]);
  fa FA_00000743 (S[606],C[603],S[607],S[743],C[743]);
  fa FA_00000744 (C[604],S[608],C[605],S[744],C[744]);
  fa FA_00000745 (S[609],C[606],S[610],S[745],C[745]);
  fa FA_00000746 (C[607],S[611],C[608],S[746],C[746]);
  fa FA_00000747 (S[612],C[609],S[613],S[747],C[747]);
  fa FA_00000748 (C[610],S[614],C[611],S[748],C[748]);
  fa FA_00000749 (S[615],C[612],S[616],S[749],C[749]);
  fa FA_00000750 (C[613],S[617],C[614],S[750],C[750]);
  fa FA_00000751 (S[618],C[615],S[619],S[751],C[751]);
  fa FA_00000752 (C[616],S[620],C[617],S[752],C[752]);
  fa FA_00000753 (S[621],C[618],S[622],S[753],C[753]);
  fa FA_00000754 (C[619],S[623],C[620],S[754],C[754]);
  fa FA_00000755 (S[624],C[621],S[625],S[755],C[755]);
  fa FA_00000756 (C[622],S[626],C[623],S[756],C[756]);
  fa FA_00000757 (S[627],C[624],S[628],S[757],C[757]);
  fa FA_00000758 (C[625],S[629],C[626],S[758],C[758]);
  fa FA_00000759 (S[630],C[627],S[631],S[759],C[759]);
  fa FA_00000760 (C[628],S[632],C[629],S[760],C[760]);
  fa FA_00000761 (S[633],C[630],S[634],S[761],C[761]);
  fa FA_00000762 (C[631],S[635],C[632],S[762],C[762]);
  fa FA_00000763 (S[636],C[633],S[637],S[763],C[763]);
  fa FA_00000764 (C[634],S[638],C[635],S[764],C[764]);
  fa FA_00000765 (S[639],C[636],S[640],S[765],C[765]);
  fa FA_00000766 (C[637],S[641],C[638],S[766],C[766]);
  fa FA_00000767 (S[642],C[639],S[643],S[767],C[767]);
  fa FA_00000768 (C[640],S[644],C[641],S[768],C[768]);
  fa FA_00000769 (S[645],C[642],S[646],S[769],C[769]);
  fa FA_00000770 (C[643],S[647],C[644],S[770],C[770]);
  fa FA_00000771 (S[648],C[645],S[649],S[771],C[771]);
  fa FA_00000772 (C[646],S[650],C[647],S[772],C[772]);
  fa FA_00000773 (S[651],C[648],S[652],S[773],C[773]);
  fa FA_00000774 (C[649],S[653],C[650],S[774],C[774]);
  fa FA_00000775 (S[654],C[651],S[655],S[775],C[775]);
  fa FA_00000776 (C[652],S[656],C[653],S[776],C[776]);
  fa FA_00000777 (S[657],C[654],S[658],S[777],C[777]);
  fa FA_00000778 (C[655],S[659],C[656],S[778],C[778]);
  fa FA_00000779 (S[660],C[657],S[661],S[779],C[779]);
  fa FA_00000780 (C[658],S[662],C[659],S[780],C[780]);
  fa FA_00000781 (S[663],C[660],S[664],S[781],C[781]);
  fa FA_00000782 (C[661],S[665],C[662],S[782],C[782]);
  fa FA_00000783 (S[666],C[663],S[667],S[783],C[783]);
  fa FA_00000784 (C[664],S[668],C[665],S[784],C[784]);
  fa FA_00000785 (S[669],C[666],S[670],S[785],C[785]);
  fa FA_00000786 (C[667],S[671],C[668],S[786],C[786]);
  fa FA_00000787 (S[672],C[669],S[673],S[787],C[787]);
  fa FA_00000788 (C[670],S[674],C[671],S[788],C[788]);
  fa FA_00000789 (S[675],C[672],S[676],S[789],C[789]);
  fa FA_00000790 (C[673],S[677],C[674],S[790],C[790]);
  fa FA_00000791 (S[678],C[675],S[679],S[791],C[791]);
  fa FA_00000792 (C[676],S[680],C[677],S[792],C[792]);
  fa FA_00000793 (S[681],C[678],S[682],S[793],C[793]);
  fa FA_00000794 (C[679],S[683],C[680],S[794],C[794]);
  fa FA_00000795 (S[684],C[681],S[685],S[795],C[795]);
  fa FA_00000796 (C[682],S[686],C[683],S[796],C[796]);
  fa FA_00000797 (S[687],C[684],S[688],S[797],C[797]);
  fa FA_00000798 (C[685],S[689],C[686],S[798],C[798]);
  fa FA_00000799 (S[690],C[687],S[691],S[799],C[799]);
  fa FA_00000800 (C[688],S[692],C[689],S[800],C[800]);
  fa FA_00000801 (S[693],C[690],S[694],S[801],C[801]);
  fa FA_00000802 (C[691],S[695],C[692],S[802],C[802]);
  fa FA_00000803 (S[696],C[693],S[697],S[803],C[803]);
  fa FA_00000804 (C[694],S[698],C[695],S[804],C[804]);
  fa FA_00000805 (S[699],C[696],S[700],S[805],C[805]);
  fa FA_00000806 (C[697],C[698],P[31][25],S[806],C[806]);
  fa FA_00000807 (S[701],C[699],C[700],S[807],C[807]);
  fa FA_00000808 (P[29][28],P[30][27],P[31][26],S[808],C[808]);
  fa FA_00000809 (C[701],P[27][31],P[28][30],S[809],C[809]);
  fa FA_00000810 (P[29][29],P[30][28],P[31][27],S[810],C[810]);
  fa FA_00000811 (P[28][31],P[29][30],P[30][29],S[811],C[811]);
  ha HA_00000812 (P[0][3],P[1][2],S[812],C[812]);
  fa FA_00000813 (S[702],P[2][2],P[3][1],S[813],C[813]);
  fa FA_00000814 (S[703],C[702],S[704],S[814],C[814]);
  fa FA_00000815 (S[705],C[703],S[706],S[815],C[815]);
  fa FA_00000816 (S[707],C[705],S[708],S[816],C[816]);
  fa FA_00000817 (S[709],C[707],S[710],S[817],C[817]);
  fa FA_00000818 (S[711],C[709],S[712],S[818],C[818]);
  fa FA_00000819 (S[713],C[711],S[714],S[819],C[819]);
  fa FA_00000820 (S[715],C[713],S[716],S[820],C[820]);
  fa FA_00000821 (S[717],C[715],S[718],S[821],C[821]);
  fa FA_00000822 (S[719],C[717],S[720],S[822],C[822]);
  fa FA_00000823 (S[721],C[719],S[722],S[823],C[823]);
  fa FA_00000824 (S[723],C[721],S[724],S[824],C[824]);
  fa FA_00000825 (S[725],C[723],S[726],S[825],C[825]);
  fa FA_00000826 (S[727],C[725],S[728],S[826],C[826]);
  fa FA_00000827 (S[729],C[727],S[730],S[827],C[827]);
  fa FA_00000828 (S[731],C[729],S[732],S[828],C[828]);
  fa FA_00000829 (S[733],C[731],S[734],S[829],C[829]);
  fa FA_00000830 (S[735],C[733],S[736],S[830],C[830]);
  fa FA_00000831 (S[737],C[735],S[738],S[831],C[831]);
  fa FA_00000832 (S[739],C[737],S[740],S[832],C[832]);
  fa FA_00000833 (S[741],C[739],S[742],S[833],C[833]);
  fa FA_00000834 (S[743],C[741],S[744],S[834],C[834]);
  fa FA_00000835 (S[745],C[743],S[746],S[835],C[835]);
  fa FA_00000836 (S[747],C[745],S[748],S[836],C[836]);
  fa FA_00000837 (S[749],C[747],S[750],S[837],C[837]);
  fa FA_00000838 (S[751],C[749],S[752],S[838],C[838]);
  fa FA_00000839 (S[753],C[751],S[754],S[839],C[839]);
  fa FA_00000840 (S[755],C[753],S[756],S[840],C[840]);
  fa FA_00000841 (S[757],C[755],S[758],S[841],C[841]);
  fa FA_00000842 (S[759],C[757],S[760],S[842],C[842]);
  fa FA_00000843 (S[761],C[759],S[762],S[843],C[843]);
  fa FA_00000844 (S[763],C[761],S[764],S[844],C[844]);
  fa FA_00000845 (S[765],C[763],S[766],S[845],C[845]);
  fa FA_00000846 (S[767],C[765],S[768],S[846],C[846]);
  fa FA_00000847 (S[769],C[767],S[770],S[847],C[847]);
  fa FA_00000848 (S[771],C[769],S[772],S[848],C[848]);
  fa FA_00000849 (S[773],C[771],S[774],S[849],C[849]);
  fa FA_00000850 (S[775],C[773],S[776],S[850],C[850]);
  fa FA_00000851 (S[777],C[775],S[778],S[851],C[851]);
  fa FA_00000852 (S[779],C[777],S[780],S[852],C[852]);
  fa FA_00000853 (S[781],C[779],S[782],S[853],C[853]);
  fa FA_00000854 (S[783],C[781],S[784],S[854],C[854]);
  fa FA_00000855 (S[785],C[783],S[786],S[855],C[855]);
  fa FA_00000856 (S[787],C[785],S[788],S[856],C[856]);
  fa FA_00000857 (S[789],C[787],S[790],S[857],C[857]);
  fa FA_00000858 (S[791],C[789],S[792],S[858],C[858]);
  fa FA_00000859 (S[793],C[791],S[794],S[859],C[859]);
  fa FA_00000860 (S[795],C[793],S[796],S[860],C[860]);
  fa FA_00000861 (S[797],C[795],S[798],S[861],C[861]);
  fa FA_00000862 (S[799],C[797],S[800],S[862],C[862]);
  fa FA_00000863 (S[801],C[799],S[802],S[863],C[863]);
  fa FA_00000864 (S[803],C[801],S[804],S[864],C[864]);
  fa FA_00000865 (S[805],C[803],S[806],S[865],C[865]);
  fa FA_00000866 (S[807],C[805],S[808],S[866],C[866]);
  fa FA_00000867 (S[809],C[807],S[810],S[867],C[867]);
  fa FA_00000868 (S[811],C[809],C[810],S[868],C[868]);
  fa FA_00000869 (C[811],P[29][31],P[30][30],S[869],C[869]);
  ha HA_00000870 (P[0][2],P[1][1],S[870],C[870]);
  fa FA_00000871 (S[812],P[2][1],P[3][0],S[871],C[871]);
  fa FA_00000872 (S[813],C[812],P[4][0],S[872],C[872]);
  fa FA_00000873 (S[814],C[813],P[5][0],S[873],C[873]);
  fa FA_00000874 (S[815],C[814],C[704],S[874],C[874]);
  fa FA_00000875 (S[816],C[815],C[706],S[875],C[875]);
  fa FA_00000876 (S[817],C[816],C[708],S[876],C[876]);
  fa FA_00000877 (S[818],C[817],C[710],S[877],C[877]);
  fa FA_00000878 (S[819],C[818],C[712],S[878],C[878]);
  fa FA_00000879 (S[820],C[819],C[714],S[879],C[879]);
  fa FA_00000880 (S[821],C[820],C[716],S[880],C[880]);
  fa FA_00000881 (S[822],C[821],C[718],S[881],C[881]);
  fa FA_00000882 (S[823],C[822],C[720],S[882],C[882]);
  fa FA_00000883 (S[824],C[823],C[722],S[883],C[883]);
  fa FA_00000884 (S[825],C[824],C[724],S[884],C[884]);
  fa FA_00000885 (S[826],C[825],C[726],S[885],C[885]);
  fa FA_00000886 (S[827],C[826],C[728],S[886],C[886]);
  fa FA_00000887 (S[828],C[827],C[730],S[887],C[887]);
  fa FA_00000888 (S[829],C[828],C[732],S[888],C[888]);
  fa FA_00000889 (S[830],C[829],C[734],S[889],C[889]);
  fa FA_00000890 (S[831],C[830],C[736],S[890],C[890]);
  fa FA_00000891 (S[832],C[831],C[738],S[891],C[891]);
  fa FA_00000892 (S[833],C[832],C[740],S[892],C[892]);
  fa FA_00000893 (S[834],C[833],C[742],S[893],C[893]);
  fa FA_00000894 (S[835],C[834],C[744],S[894],C[894]);
  fa FA_00000895 (S[836],C[835],C[746],S[895],C[895]);
  fa FA_00000896 (S[837],C[836],C[748],S[896],C[896]);
  fa FA_00000897 (S[838],C[837],C[750],S[897],C[897]);
  fa FA_00000898 (S[839],C[838],C[752],S[898],C[898]);
  fa FA_00000899 (S[840],C[839],C[754],S[899],C[899]);
  fa FA_00000900 (S[841],C[840],C[756],S[900],C[900]);
  fa FA_00000901 (S[842],C[841],C[758],S[901],C[901]);
  fa FA_00000902 (S[843],C[842],C[760],S[902],C[902]);
  fa FA_00000903 (S[844],C[843],C[762],S[903],C[903]);
  fa FA_00000904 (S[845],C[844],C[764],S[904],C[904]);
  fa FA_00000905 (S[846],C[845],C[766],S[905],C[905]);
  fa FA_00000906 (S[847],C[846],C[768],S[906],C[906]);
  fa FA_00000907 (S[848],C[847],C[770],S[907],C[907]);
  fa FA_00000908 (S[849],C[848],C[772],S[908],C[908]);
  fa FA_00000909 (S[850],C[849],C[774],S[909],C[909]);
  fa FA_00000910 (S[851],C[850],C[776],S[910],C[910]);
  fa FA_00000911 (S[852],C[851],C[778],S[911],C[911]);
  fa FA_00000912 (S[853],C[852],C[780],S[912],C[912]);
  fa FA_00000913 (S[854],C[853],C[782],S[913],C[913]);
  fa FA_00000914 (S[855],C[854],C[784],S[914],C[914]);
  fa FA_00000915 (S[856],C[855],C[786],S[915],C[915]);
  fa FA_00000916 (S[857],C[856],C[788],S[916],C[916]);
  fa FA_00000917 (S[858],C[857],C[790],S[917],C[917]);
  fa FA_00000918 (S[859],C[858],C[792],S[918],C[918]);
  fa FA_00000919 (S[860],C[859],C[794],S[919],C[919]);
  fa FA_00000920 (S[861],C[860],C[796],S[920],C[920]);
  fa FA_00000921 (S[862],C[861],C[798],S[921],C[921]);
  fa FA_00000922 (S[863],C[862],C[800],S[922],C[922]);
  fa FA_00000923 (S[864],C[863],C[802],S[923],C[923]);
  fa FA_00000924 (S[865],C[864],C[804],S[924],C[924]);
  fa FA_00000925 (S[866],C[865],C[806],S[925],C[925]);
  fa FA_00000926 (S[867],C[866],C[808],S[926],C[926]);
  fa FA_00000927 (S[868],C[867],P[31][28],S[927],C[927]);
  fa FA_00000928 (S[869],C[868],P[31][29],S[928],C[928]);
  fa FA_00000929 (C[869],P[30][31],P[31][30],S[929],C[929]);

  assign z0[0] = P[0][0];
  assign z0[1] = P[0][1];
  assign z0[2] = S[870];
  assign z0[3] = S[871];
  assign z0[4] = S[872];
  assign z0[5] = S[873];
  assign z0[6] = S[874];
  assign z0[7] = S[875];
  assign z0[8] = S[876];
  assign z0[9] = S[877];
  assign z0[10] = S[878];
  assign z0[11] = S[879];
  assign z0[12] = S[880];
  assign z0[13] = S[881];
  assign z0[14] = S[882];
  assign z0[15] = S[883];
  assign z0[16] = S[884];
  assign z0[17] = S[885];
  assign z0[18] = S[886];
  assign z0[19] = S[887];
  assign z0[20] = S[888];
  assign z0[21] = S[889];
  assign z0[22] = S[890];
  assign z0[23] = S[891];
  assign z0[24] = S[892];
  assign z0[25] = S[893];
  assign z0[26] = S[894];
  assign z0[27] = S[895];
  assign z0[28] = S[896];
  assign z0[29] = S[897];
  assign z0[30] = S[898];
  assign z0[31] = S[899];
  assign z0[32] = S[900];
  assign z0[33] = S[901];
  assign z0[34] = S[902];
  assign z0[35] = S[903];
  assign z0[36] = S[904];
  assign z0[37] = S[905];
  assign z0[38] = S[906];
  assign z0[39] = S[907];
  assign z0[40] = S[908];
  assign z0[41] = S[909];
  assign z0[42] = S[910];
  assign z0[43] = S[911];
  assign z0[44] = S[912];
  assign z0[45] = S[913];
  assign z0[46] = S[914];
  assign z0[47] = S[915];
  assign z0[48] = S[916];
  assign z0[49] = S[917];
  assign z0[50] = S[918];
  assign z0[51] = S[919];
  assign z0[52] = S[920];
  assign z0[53] = S[921];
  assign z0[54] = S[922];
  assign z0[55] = S[923];
  assign z0[56] = S[924];
  assign z0[57] = S[925];
  assign z0[58] = S[926];
  assign z0[59] = S[927];
  assign z0[60] = S[928];
  assign z0[61] = S[929];
  assign z0[62] = C[929];
  assign z0[63] = 0;
  assign z1[0] = 0;
  assign z1[1] = P[1][0];
  assign z1[2] = P[2][0];
  assign z1[3] = C[870];
  assign z1[4] = C[871];
  assign z1[5] = C[872];
  assign z1[6] = C[873];
  assign z1[7] = C[874];
  assign z1[8] = C[875];
  assign z1[9] = C[876];
  assign z1[10] = C[877];
  assign z1[11] = C[878];
  assign z1[12] = C[879];
  assign z1[13] = C[880];
  assign z1[14] = C[881];
  assign z1[15] = C[882];
  assign z1[16] = C[883];
  assign z1[17] = C[884];
  assign z1[18] = C[885];
  assign z1[19] = C[886];
  assign z1[20] = C[887];
  assign z1[21] = C[888];
  assign z1[22] = C[889];
  assign z1[23] = C[890];
  assign z1[24] = C[891];
  assign z1[25] = C[892];
  assign z1[26] = C[893];
  assign z1[27] = C[894];
  assign z1[28] = C[895];
  assign z1[29] = C[896];
  assign z1[30] = C[897];
  assign z1[31] = C[898];
  assign z1[32] = C[899];
  assign z1[33] = C[900];
  assign z1[34] = C[901];
  assign z1[35] = C[902];
  assign z1[36] = C[903];
  assign z1[37] = C[904];
  assign z1[38] = C[905];
  assign z1[39] = C[906];
  assign z1[40] = C[907];
  assign z1[41] = C[908];
  assign z1[42] = C[909];
  assign z1[43] = C[910];
  assign z1[44] = C[911];
  assign z1[45] = C[912];
  assign z1[46] = C[913];
  assign z1[47] = C[914];
  assign z1[48] = C[915];
  assign z1[49] = C[916];
  assign z1[50] = C[917];
  assign z1[51] = C[918];
  assign z1[52] = C[919];
  assign z1[53] = C[920];
  assign z1[54] = C[921];
  assign z1[55] = C[922];
  assign z1[56] = C[923];
  assign z1[57] = C[924];
  assign z1[58] = C[925];
  assign z1[59] = C[926];
  assign z1[60] = C[927];
  assign z1[61] = C[928];
  assign z1[62] = P[31][31];
  assign z1[63] = 0;

endmodule


module wallace
(
  input  [31 : 0] x,
  input  [31 : 0] y,
  output [63 : 0] z0,
  output [63 : 0] z1
);

  wire [31 : 0] P [0 : 31];

  wire [1061 : 0] S;
  wire [1061 : 0] C;

  assign P[0][0] = x[0] & y[0];
  assign P[0][1] = x[0] & y[1];
  assign P[0][2] = x[0] & y[2];
  assign P[0][3] = x[0] & y[3];
  assign P[0][4] = x[0] & y[4];
  assign P[0][5] = x[0] & y[5];
  assign P[0][6] = x[0] & y[6];
  assign P[0][7] = x[0] & y[7];
  assign P[0][8] = x[0] & y[8];
  assign P[0][9] = x[0] & y[9];
  assign P[0][10] = x[0] & y[10];
  assign P[0][11] = x[0] & y[11];
  assign P[0][12] = x[0] & y[12];
  assign P[0][13] = x[0] & y[13];
  assign P[0][14] = x[0] & y[14];
  assign P[0][15] = x[0] & y[15];
  assign P[0][16] = x[0] & y[16];
  assign P[0][17] = x[0] & y[17];
  assign P[0][18] = x[0] & y[18];
  assign P[0][19] = x[0] & y[19];
  assign P[0][20] = x[0] & y[20];
  assign P[0][21] = x[0] & y[21];
  assign P[0][22] = x[0] & y[22];
  assign P[0][23] = x[0] & y[23];
  assign P[0][24] = x[0] & y[24];
  assign P[0][25] = x[0] & y[25];
  assign P[0][26] = x[0] & y[26];
  assign P[0][27] = x[0] & y[27];
  assign P[0][28] = x[0] & y[28];
  assign P[0][29] = x[0] & y[29];
  assign P[0][30] = x[0] & y[30];
  assign P[0][31] = x[0] & y[31];
  assign P[1][0] = x[1] & y[0];
  assign P[1][1] = x[1] & y[1];
  assign P[1][2] = x[1] & y[2];
  assign P[1][3] = x[1] & y[3];
  assign P[1][4] = x[1] & y[4];
  assign P[1][5] = x[1] & y[5];
  assign P[1][6] = x[1] & y[6];
  assign P[1][7] = x[1] & y[7];
  assign P[1][8] = x[1] & y[8];
  assign P[1][9] = x[1] & y[9];
  assign P[1][10] = x[1] & y[10];
  assign P[1][11] = x[1] & y[11];
  assign P[1][12] = x[1] & y[12];
  assign P[1][13] = x[1] & y[13];
  assign P[1][14] = x[1] & y[14];
  assign P[1][15] = x[1] & y[15];
  assign P[1][16] = x[1] & y[16];
  assign P[1][17] = x[1] & y[17];
  assign P[1][18] = x[1] & y[18];
  assign P[1][19] = x[1] & y[19];
  assign P[1][20] = x[1] & y[20];
  assign P[1][21] = x[1] & y[21];
  assign P[1][22] = x[1] & y[22];
  assign P[1][23] = x[1] & y[23];
  assign P[1][24] = x[1] & y[24];
  assign P[1][25] = x[1] & y[25];
  assign P[1][26] = x[1] & y[26];
  assign P[1][27] = x[1] & y[27];
  assign P[1][28] = x[1] & y[28];
  assign P[1][29] = x[1] & y[29];
  assign P[1][30] = x[1] & y[30];
  assign P[1][31] = x[1] & y[31];
  assign P[2][0] = x[2] & y[0];
  assign P[2][1] = x[2] & y[1];
  assign P[2][2] = x[2] & y[2];
  assign P[2][3] = x[2] & y[3];
  assign P[2][4] = x[2] & y[4];
  assign P[2][5] = x[2] & y[5];
  assign P[2][6] = x[2] & y[6];
  assign P[2][7] = x[2] & y[7];
  assign P[2][8] = x[2] & y[8];
  assign P[2][9] = x[2] & y[9];
  assign P[2][10] = x[2] & y[10];
  assign P[2][11] = x[2] & y[11];
  assign P[2][12] = x[2] & y[12];
  assign P[2][13] = x[2] & y[13];
  assign P[2][14] = x[2] & y[14];
  assign P[2][15] = x[2] & y[15];
  assign P[2][16] = x[2] & y[16];
  assign P[2][17] = x[2] & y[17];
  assign P[2][18] = x[2] & y[18];
  assign P[2][19] = x[2] & y[19];
  assign P[2][20] = x[2] & y[20];
  assign P[2][21] = x[2] & y[21];
  assign P[2][22] = x[2] & y[22];
  assign P[2][23] = x[2] & y[23];
  assign P[2][24] = x[2] & y[24];
  assign P[2][25] = x[2] & y[25];
  assign P[2][26] = x[2] & y[26];
  assign P[2][27] = x[2] & y[27];
  assign P[2][28] = x[2] & y[28];
  assign P[2][29] = x[2] & y[29];
  assign P[2][30] = x[2] & y[30];
  assign P[2][31] = x[2] & y[31];
  assign P[3][0] = x[3] & y[0];
  assign P[3][1] = x[3] & y[1];
  assign P[3][2] = x[3] & y[2];
  assign P[3][3] = x[3] & y[3];
  assign P[3][4] = x[3] & y[4];
  assign P[3][5] = x[3] & y[5];
  assign P[3][6] = x[3] & y[6];
  assign P[3][7] = x[3] & y[7];
  assign P[3][8] = x[3] & y[8];
  assign P[3][9] = x[3] & y[9];
  assign P[3][10] = x[3] & y[10];
  assign P[3][11] = x[3] & y[11];
  assign P[3][12] = x[3] & y[12];
  assign P[3][13] = x[3] & y[13];
  assign P[3][14] = x[3] & y[14];
  assign P[3][15] = x[3] & y[15];
  assign P[3][16] = x[3] & y[16];
  assign P[3][17] = x[3] & y[17];
  assign P[3][18] = x[3] & y[18];
  assign P[3][19] = x[3] & y[19];
  assign P[3][20] = x[3] & y[20];
  assign P[3][21] = x[3] & y[21];
  assign P[3][22] = x[3] & y[22];
  assign P[3][23] = x[3] & y[23];
  assign P[3][24] = x[3] & y[24];
  assign P[3][25] = x[3] & y[25];
  assign P[3][26] = x[3] & y[26];
  assign P[3][27] = x[3] & y[27];
  assign P[3][28] = x[3] & y[28];
  assign P[3][29] = x[3] & y[29];
  assign P[3][30] = x[3] & y[30];
  assign P[3][31] = x[3] & y[31];
  assign P[4][0] = x[4] & y[0];
  assign P[4][1] = x[4] & y[1];
  assign P[4][2] = x[4] & y[2];
  assign P[4][3] = x[4] & y[3];
  assign P[4][4] = x[4] & y[4];
  assign P[4][5] = x[4] & y[5];
  assign P[4][6] = x[4] & y[6];
  assign P[4][7] = x[4] & y[7];
  assign P[4][8] = x[4] & y[8];
  assign P[4][9] = x[4] & y[9];
  assign P[4][10] = x[4] & y[10];
  assign P[4][11] = x[4] & y[11];
  assign P[4][12] = x[4] & y[12];
  assign P[4][13] = x[4] & y[13];
  assign P[4][14] = x[4] & y[14];
  assign P[4][15] = x[4] & y[15];
  assign P[4][16] = x[4] & y[16];
  assign P[4][17] = x[4] & y[17];
  assign P[4][18] = x[4] & y[18];
  assign P[4][19] = x[4] & y[19];
  assign P[4][20] = x[4] & y[20];
  assign P[4][21] = x[4] & y[21];
  assign P[4][22] = x[4] & y[22];
  assign P[4][23] = x[4] & y[23];
  assign P[4][24] = x[4] & y[24];
  assign P[4][25] = x[4] & y[25];
  assign P[4][26] = x[4] & y[26];
  assign P[4][27] = x[4] & y[27];
  assign P[4][28] = x[4] & y[28];
  assign P[4][29] = x[4] & y[29];
  assign P[4][30] = x[4] & y[30];
  assign P[4][31] = x[4] & y[31];
  assign P[5][0] = x[5] & y[0];
  assign P[5][1] = x[5] & y[1];
  assign P[5][2] = x[5] & y[2];
  assign P[5][3] = x[5] & y[3];
  assign P[5][4] = x[5] & y[4];
  assign P[5][5] = x[5] & y[5];
  assign P[5][6] = x[5] & y[6];
  assign P[5][7] = x[5] & y[7];
  assign P[5][8] = x[5] & y[8];
  assign P[5][9] = x[5] & y[9];
  assign P[5][10] = x[5] & y[10];
  assign P[5][11] = x[5] & y[11];
  assign P[5][12] = x[5] & y[12];
  assign P[5][13] = x[5] & y[13];
  assign P[5][14] = x[5] & y[14];
  assign P[5][15] = x[5] & y[15];
  assign P[5][16] = x[5] & y[16];
  assign P[5][17] = x[5] & y[17];
  assign P[5][18] = x[5] & y[18];
  assign P[5][19] = x[5] & y[19];
  assign P[5][20] = x[5] & y[20];
  assign P[5][21] = x[5] & y[21];
  assign P[5][22] = x[5] & y[22];
  assign P[5][23] = x[5] & y[23];
  assign P[5][24] = x[5] & y[24];
  assign P[5][25] = x[5] & y[25];
  assign P[5][26] = x[5] & y[26];
  assign P[5][27] = x[5] & y[27];
  assign P[5][28] = x[5] & y[28];
  assign P[5][29] = x[5] & y[29];
  assign P[5][30] = x[5] & y[30];
  assign P[5][31] = x[5] & y[31];
  assign P[6][0] = x[6] & y[0];
  assign P[6][1] = x[6] & y[1];
  assign P[6][2] = x[6] & y[2];
  assign P[6][3] = x[6] & y[3];
  assign P[6][4] = x[6] & y[4];
  assign P[6][5] = x[6] & y[5];
  assign P[6][6] = x[6] & y[6];
  assign P[6][7] = x[6] & y[7];
  assign P[6][8] = x[6] & y[8];
  assign P[6][9] = x[6] & y[9];
  assign P[6][10] = x[6] & y[10];
  assign P[6][11] = x[6] & y[11];
  assign P[6][12] = x[6] & y[12];
  assign P[6][13] = x[6] & y[13];
  assign P[6][14] = x[6] & y[14];
  assign P[6][15] = x[6] & y[15];
  assign P[6][16] = x[6] & y[16];
  assign P[6][17] = x[6] & y[17];
  assign P[6][18] = x[6] & y[18];
  assign P[6][19] = x[6] & y[19];
  assign P[6][20] = x[6] & y[20];
  assign P[6][21] = x[6] & y[21];
  assign P[6][22] = x[6] & y[22];
  assign P[6][23] = x[6] & y[23];
  assign P[6][24] = x[6] & y[24];
  assign P[6][25] = x[6] & y[25];
  assign P[6][26] = x[6] & y[26];
  assign P[6][27] = x[6] & y[27];
  assign P[6][28] = x[6] & y[28];
  assign P[6][29] = x[6] & y[29];
  assign P[6][30] = x[6] & y[30];
  assign P[6][31] = x[6] & y[31];
  assign P[7][0] = x[7] & y[0];
  assign P[7][1] = x[7] & y[1];
  assign P[7][2] = x[7] & y[2];
  assign P[7][3] = x[7] & y[3];
  assign P[7][4] = x[7] & y[4];
  assign P[7][5] = x[7] & y[5];
  assign P[7][6] = x[7] & y[6];
  assign P[7][7] = x[7] & y[7];
  assign P[7][8] = x[7] & y[8];
  assign P[7][9] = x[7] & y[9];
  assign P[7][10] = x[7] & y[10];
  assign P[7][11] = x[7] & y[11];
  assign P[7][12] = x[7] & y[12];
  assign P[7][13] = x[7] & y[13];
  assign P[7][14] = x[7] & y[14];
  assign P[7][15] = x[7] & y[15];
  assign P[7][16] = x[7] & y[16];
  assign P[7][17] = x[7] & y[17];
  assign P[7][18] = x[7] & y[18];
  assign P[7][19] = x[7] & y[19];
  assign P[7][20] = x[7] & y[20];
  assign P[7][21] = x[7] & y[21];
  assign P[7][22] = x[7] & y[22];
  assign P[7][23] = x[7] & y[23];
  assign P[7][24] = x[7] & y[24];
  assign P[7][25] = x[7] & y[25];
  assign P[7][26] = x[7] & y[26];
  assign P[7][27] = x[7] & y[27];
  assign P[7][28] = x[7] & y[28];
  assign P[7][29] = x[7] & y[29];
  assign P[7][30] = x[7] & y[30];
  assign P[7][31] = x[7] & y[31];
  assign P[8][0] = x[8] & y[0];
  assign P[8][1] = x[8] & y[1];
  assign P[8][2] = x[8] & y[2];
  assign P[8][3] = x[8] & y[3];
  assign P[8][4] = x[8] & y[4];
  assign P[8][5] = x[8] & y[5];
  assign P[8][6] = x[8] & y[6];
  assign P[8][7] = x[8] & y[7];
  assign P[8][8] = x[8] & y[8];
  assign P[8][9] = x[8] & y[9];
  assign P[8][10] = x[8] & y[10];
  assign P[8][11] = x[8] & y[11];
  assign P[8][12] = x[8] & y[12];
  assign P[8][13] = x[8] & y[13];
  assign P[8][14] = x[8] & y[14];
  assign P[8][15] = x[8] & y[15];
  assign P[8][16] = x[8] & y[16];
  assign P[8][17] = x[8] & y[17];
  assign P[8][18] = x[8] & y[18];
  assign P[8][19] = x[8] & y[19];
  assign P[8][20] = x[8] & y[20];
  assign P[8][21] = x[8] & y[21];
  assign P[8][22] = x[8] & y[22];
  assign P[8][23] = x[8] & y[23];
  assign P[8][24] = x[8] & y[24];
  assign P[8][25] = x[8] & y[25];
  assign P[8][26] = x[8] & y[26];
  assign P[8][27] = x[8] & y[27];
  assign P[8][28] = x[8] & y[28];
  assign P[8][29] = x[8] & y[29];
  assign P[8][30] = x[8] & y[30];
  assign P[8][31] = x[8] & y[31];
  assign P[9][0] = x[9] & y[0];
  assign P[9][1] = x[9] & y[1];
  assign P[9][2] = x[9] & y[2];
  assign P[9][3] = x[9] & y[3];
  assign P[9][4] = x[9] & y[4];
  assign P[9][5] = x[9] & y[5];
  assign P[9][6] = x[9] & y[6];
  assign P[9][7] = x[9] & y[7];
  assign P[9][8] = x[9] & y[8];
  assign P[9][9] = x[9] & y[9];
  assign P[9][10] = x[9] & y[10];
  assign P[9][11] = x[9] & y[11];
  assign P[9][12] = x[9] & y[12];
  assign P[9][13] = x[9] & y[13];
  assign P[9][14] = x[9] & y[14];
  assign P[9][15] = x[9] & y[15];
  assign P[9][16] = x[9] & y[16];
  assign P[9][17] = x[9] & y[17];
  assign P[9][18] = x[9] & y[18];
  assign P[9][19] = x[9] & y[19];
  assign P[9][20] = x[9] & y[20];
  assign P[9][21] = x[9] & y[21];
  assign P[9][22] = x[9] & y[22];
  assign P[9][23] = x[9] & y[23];
  assign P[9][24] = x[9] & y[24];
  assign P[9][25] = x[9] & y[25];
  assign P[9][26] = x[9] & y[26];
  assign P[9][27] = x[9] & y[27];
  assign P[9][28] = x[9] & y[28];
  assign P[9][29] = x[9] & y[29];
  assign P[9][30] = x[9] & y[30];
  assign P[9][31] = x[9] & y[31];
  assign P[10][0] = x[10] & y[0];
  assign P[10][1] = x[10] & y[1];
  assign P[10][2] = x[10] & y[2];
  assign P[10][3] = x[10] & y[3];
  assign P[10][4] = x[10] & y[4];
  assign P[10][5] = x[10] & y[5];
  assign P[10][6] = x[10] & y[6];
  assign P[10][7] = x[10] & y[7];
  assign P[10][8] = x[10] & y[8];
  assign P[10][9] = x[10] & y[9];
  assign P[10][10] = x[10] & y[10];
  assign P[10][11] = x[10] & y[11];
  assign P[10][12] = x[10] & y[12];
  assign P[10][13] = x[10] & y[13];
  assign P[10][14] = x[10] & y[14];
  assign P[10][15] = x[10] & y[15];
  assign P[10][16] = x[10] & y[16];
  assign P[10][17] = x[10] & y[17];
  assign P[10][18] = x[10] & y[18];
  assign P[10][19] = x[10] & y[19];
  assign P[10][20] = x[10] & y[20];
  assign P[10][21] = x[10] & y[21];
  assign P[10][22] = x[10] & y[22];
  assign P[10][23] = x[10] & y[23];
  assign P[10][24] = x[10] & y[24];
  assign P[10][25] = x[10] & y[25];
  assign P[10][26] = x[10] & y[26];
  assign P[10][27] = x[10] & y[27];
  assign P[10][28] = x[10] & y[28];
  assign P[10][29] = x[10] & y[29];
  assign P[10][30] = x[10] & y[30];
  assign P[10][31] = x[10] & y[31];
  assign P[11][0] = x[11] & y[0];
  assign P[11][1] = x[11] & y[1];
  assign P[11][2] = x[11] & y[2];
  assign P[11][3] = x[11] & y[3];
  assign P[11][4] = x[11] & y[4];
  assign P[11][5] = x[11] & y[5];
  assign P[11][6] = x[11] & y[6];
  assign P[11][7] = x[11] & y[7];
  assign P[11][8] = x[11] & y[8];
  assign P[11][9] = x[11] & y[9];
  assign P[11][10] = x[11] & y[10];
  assign P[11][11] = x[11] & y[11];
  assign P[11][12] = x[11] & y[12];
  assign P[11][13] = x[11] & y[13];
  assign P[11][14] = x[11] & y[14];
  assign P[11][15] = x[11] & y[15];
  assign P[11][16] = x[11] & y[16];
  assign P[11][17] = x[11] & y[17];
  assign P[11][18] = x[11] & y[18];
  assign P[11][19] = x[11] & y[19];
  assign P[11][20] = x[11] & y[20];
  assign P[11][21] = x[11] & y[21];
  assign P[11][22] = x[11] & y[22];
  assign P[11][23] = x[11] & y[23];
  assign P[11][24] = x[11] & y[24];
  assign P[11][25] = x[11] & y[25];
  assign P[11][26] = x[11] & y[26];
  assign P[11][27] = x[11] & y[27];
  assign P[11][28] = x[11] & y[28];
  assign P[11][29] = x[11] & y[29];
  assign P[11][30] = x[11] & y[30];
  assign P[11][31] = x[11] & y[31];
  assign P[12][0] = x[12] & y[0];
  assign P[12][1] = x[12] & y[1];
  assign P[12][2] = x[12] & y[2];
  assign P[12][3] = x[12] & y[3];
  assign P[12][4] = x[12] & y[4];
  assign P[12][5] = x[12] & y[5];
  assign P[12][6] = x[12] & y[6];
  assign P[12][7] = x[12] & y[7];
  assign P[12][8] = x[12] & y[8];
  assign P[12][9] = x[12] & y[9];
  assign P[12][10] = x[12] & y[10];
  assign P[12][11] = x[12] & y[11];
  assign P[12][12] = x[12] & y[12];
  assign P[12][13] = x[12] & y[13];
  assign P[12][14] = x[12] & y[14];
  assign P[12][15] = x[12] & y[15];
  assign P[12][16] = x[12] & y[16];
  assign P[12][17] = x[12] & y[17];
  assign P[12][18] = x[12] & y[18];
  assign P[12][19] = x[12] & y[19];
  assign P[12][20] = x[12] & y[20];
  assign P[12][21] = x[12] & y[21];
  assign P[12][22] = x[12] & y[22];
  assign P[12][23] = x[12] & y[23];
  assign P[12][24] = x[12] & y[24];
  assign P[12][25] = x[12] & y[25];
  assign P[12][26] = x[12] & y[26];
  assign P[12][27] = x[12] & y[27];
  assign P[12][28] = x[12] & y[28];
  assign P[12][29] = x[12] & y[29];
  assign P[12][30] = x[12] & y[30];
  assign P[12][31] = x[12] & y[31];
  assign P[13][0] = x[13] & y[0];
  assign P[13][1] = x[13] & y[1];
  assign P[13][2] = x[13] & y[2];
  assign P[13][3] = x[13] & y[3];
  assign P[13][4] = x[13] & y[4];
  assign P[13][5] = x[13] & y[5];
  assign P[13][6] = x[13] & y[6];
  assign P[13][7] = x[13] & y[7];
  assign P[13][8] = x[13] & y[8];
  assign P[13][9] = x[13] & y[9];
  assign P[13][10] = x[13] & y[10];
  assign P[13][11] = x[13] & y[11];
  assign P[13][12] = x[13] & y[12];
  assign P[13][13] = x[13] & y[13];
  assign P[13][14] = x[13] & y[14];
  assign P[13][15] = x[13] & y[15];
  assign P[13][16] = x[13] & y[16];
  assign P[13][17] = x[13] & y[17];
  assign P[13][18] = x[13] & y[18];
  assign P[13][19] = x[13] & y[19];
  assign P[13][20] = x[13] & y[20];
  assign P[13][21] = x[13] & y[21];
  assign P[13][22] = x[13] & y[22];
  assign P[13][23] = x[13] & y[23];
  assign P[13][24] = x[13] & y[24];
  assign P[13][25] = x[13] & y[25];
  assign P[13][26] = x[13] & y[26];
  assign P[13][27] = x[13] & y[27];
  assign P[13][28] = x[13] & y[28];
  assign P[13][29] = x[13] & y[29];
  assign P[13][30] = x[13] & y[30];
  assign P[13][31] = x[13] & y[31];
  assign P[14][0] = x[14] & y[0];
  assign P[14][1] = x[14] & y[1];
  assign P[14][2] = x[14] & y[2];
  assign P[14][3] = x[14] & y[3];
  assign P[14][4] = x[14] & y[4];
  assign P[14][5] = x[14] & y[5];
  assign P[14][6] = x[14] & y[6];
  assign P[14][7] = x[14] & y[7];
  assign P[14][8] = x[14] & y[8];
  assign P[14][9] = x[14] & y[9];
  assign P[14][10] = x[14] & y[10];
  assign P[14][11] = x[14] & y[11];
  assign P[14][12] = x[14] & y[12];
  assign P[14][13] = x[14] & y[13];
  assign P[14][14] = x[14] & y[14];
  assign P[14][15] = x[14] & y[15];
  assign P[14][16] = x[14] & y[16];
  assign P[14][17] = x[14] & y[17];
  assign P[14][18] = x[14] & y[18];
  assign P[14][19] = x[14] & y[19];
  assign P[14][20] = x[14] & y[20];
  assign P[14][21] = x[14] & y[21];
  assign P[14][22] = x[14] & y[22];
  assign P[14][23] = x[14] & y[23];
  assign P[14][24] = x[14] & y[24];
  assign P[14][25] = x[14] & y[25];
  assign P[14][26] = x[14] & y[26];
  assign P[14][27] = x[14] & y[27];
  assign P[14][28] = x[14] & y[28];
  assign P[14][29] = x[14] & y[29];
  assign P[14][30] = x[14] & y[30];
  assign P[14][31] = x[14] & y[31];
  assign P[15][0] = x[15] & y[0];
  assign P[15][1] = x[15] & y[1];
  assign P[15][2] = x[15] & y[2];
  assign P[15][3] = x[15] & y[3];
  assign P[15][4] = x[15] & y[4];
  assign P[15][5] = x[15] & y[5];
  assign P[15][6] = x[15] & y[6];
  assign P[15][7] = x[15] & y[7];
  assign P[15][8] = x[15] & y[8];
  assign P[15][9] = x[15] & y[9];
  assign P[15][10] = x[15] & y[10];
  assign P[15][11] = x[15] & y[11];
  assign P[15][12] = x[15] & y[12];
  assign P[15][13] = x[15] & y[13];
  assign P[15][14] = x[15] & y[14];
  assign P[15][15] = x[15] & y[15];
  assign P[15][16] = x[15] & y[16];
  assign P[15][17] = x[15] & y[17];
  assign P[15][18] = x[15] & y[18];
  assign P[15][19] = x[15] & y[19];
  assign P[15][20] = x[15] & y[20];
  assign P[15][21] = x[15] & y[21];
  assign P[15][22] = x[15] & y[22];
  assign P[15][23] = x[15] & y[23];
  assign P[15][24] = x[15] & y[24];
  assign P[15][25] = x[15] & y[25];
  assign P[15][26] = x[15] & y[26];
  assign P[15][27] = x[15] & y[27];
  assign P[15][28] = x[15] & y[28];
  assign P[15][29] = x[15] & y[29];
  assign P[15][30] = x[15] & y[30];
  assign P[15][31] = x[15] & y[31];
  assign P[16][0] = x[16] & y[0];
  assign P[16][1] = x[16] & y[1];
  assign P[16][2] = x[16] & y[2];
  assign P[16][3] = x[16] & y[3];
  assign P[16][4] = x[16] & y[4];
  assign P[16][5] = x[16] & y[5];
  assign P[16][6] = x[16] & y[6];
  assign P[16][7] = x[16] & y[7];
  assign P[16][8] = x[16] & y[8];
  assign P[16][9] = x[16] & y[9];
  assign P[16][10] = x[16] & y[10];
  assign P[16][11] = x[16] & y[11];
  assign P[16][12] = x[16] & y[12];
  assign P[16][13] = x[16] & y[13];
  assign P[16][14] = x[16] & y[14];
  assign P[16][15] = x[16] & y[15];
  assign P[16][16] = x[16] & y[16];
  assign P[16][17] = x[16] & y[17];
  assign P[16][18] = x[16] & y[18];
  assign P[16][19] = x[16] & y[19];
  assign P[16][20] = x[16] & y[20];
  assign P[16][21] = x[16] & y[21];
  assign P[16][22] = x[16] & y[22];
  assign P[16][23] = x[16] & y[23];
  assign P[16][24] = x[16] & y[24];
  assign P[16][25] = x[16] & y[25];
  assign P[16][26] = x[16] & y[26];
  assign P[16][27] = x[16] & y[27];
  assign P[16][28] = x[16] & y[28];
  assign P[16][29] = x[16] & y[29];
  assign P[16][30] = x[16] & y[30];
  assign P[16][31] = x[16] & y[31];
  assign P[17][0] = x[17] & y[0];
  assign P[17][1] = x[17] & y[1];
  assign P[17][2] = x[17] & y[2];
  assign P[17][3] = x[17] & y[3];
  assign P[17][4] = x[17] & y[4];
  assign P[17][5] = x[17] & y[5];
  assign P[17][6] = x[17] & y[6];
  assign P[17][7] = x[17] & y[7];
  assign P[17][8] = x[17] & y[8];
  assign P[17][9] = x[17] & y[9];
  assign P[17][10] = x[17] & y[10];
  assign P[17][11] = x[17] & y[11];
  assign P[17][12] = x[17] & y[12];
  assign P[17][13] = x[17] & y[13];
  assign P[17][14] = x[17] & y[14];
  assign P[17][15] = x[17] & y[15];
  assign P[17][16] = x[17] & y[16];
  assign P[17][17] = x[17] & y[17];
  assign P[17][18] = x[17] & y[18];
  assign P[17][19] = x[17] & y[19];
  assign P[17][20] = x[17] & y[20];
  assign P[17][21] = x[17] & y[21];
  assign P[17][22] = x[17] & y[22];
  assign P[17][23] = x[17] & y[23];
  assign P[17][24] = x[17] & y[24];
  assign P[17][25] = x[17] & y[25];
  assign P[17][26] = x[17] & y[26];
  assign P[17][27] = x[17] & y[27];
  assign P[17][28] = x[17] & y[28];
  assign P[17][29] = x[17] & y[29];
  assign P[17][30] = x[17] & y[30];
  assign P[17][31] = x[17] & y[31];
  assign P[18][0] = x[18] & y[0];
  assign P[18][1] = x[18] & y[1];
  assign P[18][2] = x[18] & y[2];
  assign P[18][3] = x[18] & y[3];
  assign P[18][4] = x[18] & y[4];
  assign P[18][5] = x[18] & y[5];
  assign P[18][6] = x[18] & y[6];
  assign P[18][7] = x[18] & y[7];
  assign P[18][8] = x[18] & y[8];
  assign P[18][9] = x[18] & y[9];
  assign P[18][10] = x[18] & y[10];
  assign P[18][11] = x[18] & y[11];
  assign P[18][12] = x[18] & y[12];
  assign P[18][13] = x[18] & y[13];
  assign P[18][14] = x[18] & y[14];
  assign P[18][15] = x[18] & y[15];
  assign P[18][16] = x[18] & y[16];
  assign P[18][17] = x[18] & y[17];
  assign P[18][18] = x[18] & y[18];
  assign P[18][19] = x[18] & y[19];
  assign P[18][20] = x[18] & y[20];
  assign P[18][21] = x[18] & y[21];
  assign P[18][22] = x[18] & y[22];
  assign P[18][23] = x[18] & y[23];
  assign P[18][24] = x[18] & y[24];
  assign P[18][25] = x[18] & y[25];
  assign P[18][26] = x[18] & y[26];
  assign P[18][27] = x[18] & y[27];
  assign P[18][28] = x[18] & y[28];
  assign P[18][29] = x[18] & y[29];
  assign P[18][30] = x[18] & y[30];
  assign P[18][31] = x[18] & y[31];
  assign P[19][0] = x[19] & y[0];
  assign P[19][1] = x[19] & y[1];
  assign P[19][2] = x[19] & y[2];
  assign P[19][3] = x[19] & y[3];
  assign P[19][4] = x[19] & y[4];
  assign P[19][5] = x[19] & y[5];
  assign P[19][6] = x[19] & y[6];
  assign P[19][7] = x[19] & y[7];
  assign P[19][8] = x[19] & y[8];
  assign P[19][9] = x[19] & y[9];
  assign P[19][10] = x[19] & y[10];
  assign P[19][11] = x[19] & y[11];
  assign P[19][12] = x[19] & y[12];
  assign P[19][13] = x[19] & y[13];
  assign P[19][14] = x[19] & y[14];
  assign P[19][15] = x[19] & y[15];
  assign P[19][16] = x[19] & y[16];
  assign P[19][17] = x[19] & y[17];
  assign P[19][18] = x[19] & y[18];
  assign P[19][19] = x[19] & y[19];
  assign P[19][20] = x[19] & y[20];
  assign P[19][21] = x[19] & y[21];
  assign P[19][22] = x[19] & y[22];
  assign P[19][23] = x[19] & y[23];
  assign P[19][24] = x[19] & y[24];
  assign P[19][25] = x[19] & y[25];
  assign P[19][26] = x[19] & y[26];
  assign P[19][27] = x[19] & y[27];
  assign P[19][28] = x[19] & y[28];
  assign P[19][29] = x[19] & y[29];
  assign P[19][30] = x[19] & y[30];
  assign P[19][31] = x[19] & y[31];
  assign P[20][0] = x[20] & y[0];
  assign P[20][1] = x[20] & y[1];
  assign P[20][2] = x[20] & y[2];
  assign P[20][3] = x[20] & y[3];
  assign P[20][4] = x[20] & y[4];
  assign P[20][5] = x[20] & y[5];
  assign P[20][6] = x[20] & y[6];
  assign P[20][7] = x[20] & y[7];
  assign P[20][8] = x[20] & y[8];
  assign P[20][9] = x[20] & y[9];
  assign P[20][10] = x[20] & y[10];
  assign P[20][11] = x[20] & y[11];
  assign P[20][12] = x[20] & y[12];
  assign P[20][13] = x[20] & y[13];
  assign P[20][14] = x[20] & y[14];
  assign P[20][15] = x[20] & y[15];
  assign P[20][16] = x[20] & y[16];
  assign P[20][17] = x[20] & y[17];
  assign P[20][18] = x[20] & y[18];
  assign P[20][19] = x[20] & y[19];
  assign P[20][20] = x[20] & y[20];
  assign P[20][21] = x[20] & y[21];
  assign P[20][22] = x[20] & y[22];
  assign P[20][23] = x[20] & y[23];
  assign P[20][24] = x[20] & y[24];
  assign P[20][25] = x[20] & y[25];
  assign P[20][26] = x[20] & y[26];
  assign P[20][27] = x[20] & y[27];
  assign P[20][28] = x[20] & y[28];
  assign P[20][29] = x[20] & y[29];
  assign P[20][30] = x[20] & y[30];
  assign P[20][31] = x[20] & y[31];
  assign P[21][0] = x[21] & y[0];
  assign P[21][1] = x[21] & y[1];
  assign P[21][2] = x[21] & y[2];
  assign P[21][3] = x[21] & y[3];
  assign P[21][4] = x[21] & y[4];
  assign P[21][5] = x[21] & y[5];
  assign P[21][6] = x[21] & y[6];
  assign P[21][7] = x[21] & y[7];
  assign P[21][8] = x[21] & y[8];
  assign P[21][9] = x[21] & y[9];
  assign P[21][10] = x[21] & y[10];
  assign P[21][11] = x[21] & y[11];
  assign P[21][12] = x[21] & y[12];
  assign P[21][13] = x[21] & y[13];
  assign P[21][14] = x[21] & y[14];
  assign P[21][15] = x[21] & y[15];
  assign P[21][16] = x[21] & y[16];
  assign P[21][17] = x[21] & y[17];
  assign P[21][18] = x[21] & y[18];
  assign P[21][19] = x[21] & y[19];
  assign P[21][20] = x[21] & y[20];
  assign P[21][21] = x[21] & y[21];
  assign P[21][22] = x[21] & y[22];
  assign P[21][23] = x[21] & y[23];
  assign P[21][24] = x[21] & y[24];
  assign P[21][25] = x[21] & y[25];
  assign P[21][26] = x[21] & y[26];
  assign P[21][27] = x[21] & y[27];
  assign P[21][28] = x[21] & y[28];
  assign P[21][29] = x[21] & y[29];
  assign P[21][30] = x[21] & y[30];
  assign P[21][31] = x[21] & y[31];
  assign P[22][0] = x[22] & y[0];
  assign P[22][1] = x[22] & y[1];
  assign P[22][2] = x[22] & y[2];
  assign P[22][3] = x[22] & y[3];
  assign P[22][4] = x[22] & y[4];
  assign P[22][5] = x[22] & y[5];
  assign P[22][6] = x[22] & y[6];
  assign P[22][7] = x[22] & y[7];
  assign P[22][8] = x[22] & y[8];
  assign P[22][9] = x[22] & y[9];
  assign P[22][10] = x[22] & y[10];
  assign P[22][11] = x[22] & y[11];
  assign P[22][12] = x[22] & y[12];
  assign P[22][13] = x[22] & y[13];
  assign P[22][14] = x[22] & y[14];
  assign P[22][15] = x[22] & y[15];
  assign P[22][16] = x[22] & y[16];
  assign P[22][17] = x[22] & y[17];
  assign P[22][18] = x[22] & y[18];
  assign P[22][19] = x[22] & y[19];
  assign P[22][20] = x[22] & y[20];
  assign P[22][21] = x[22] & y[21];
  assign P[22][22] = x[22] & y[22];
  assign P[22][23] = x[22] & y[23];
  assign P[22][24] = x[22] & y[24];
  assign P[22][25] = x[22] & y[25];
  assign P[22][26] = x[22] & y[26];
  assign P[22][27] = x[22] & y[27];
  assign P[22][28] = x[22] & y[28];
  assign P[22][29] = x[22] & y[29];
  assign P[22][30] = x[22] & y[30];
  assign P[22][31] = x[22] & y[31];
  assign P[23][0] = x[23] & y[0];
  assign P[23][1] = x[23] & y[1];
  assign P[23][2] = x[23] & y[2];
  assign P[23][3] = x[23] & y[3];
  assign P[23][4] = x[23] & y[4];
  assign P[23][5] = x[23] & y[5];
  assign P[23][6] = x[23] & y[6];
  assign P[23][7] = x[23] & y[7];
  assign P[23][8] = x[23] & y[8];
  assign P[23][9] = x[23] & y[9];
  assign P[23][10] = x[23] & y[10];
  assign P[23][11] = x[23] & y[11];
  assign P[23][12] = x[23] & y[12];
  assign P[23][13] = x[23] & y[13];
  assign P[23][14] = x[23] & y[14];
  assign P[23][15] = x[23] & y[15];
  assign P[23][16] = x[23] & y[16];
  assign P[23][17] = x[23] & y[17];
  assign P[23][18] = x[23] & y[18];
  assign P[23][19] = x[23] & y[19];
  assign P[23][20] = x[23] & y[20];
  assign P[23][21] = x[23] & y[21];
  assign P[23][22] = x[23] & y[22];
  assign P[23][23] = x[23] & y[23];
  assign P[23][24] = x[23] & y[24];
  assign P[23][25] = x[23] & y[25];
  assign P[23][26] = x[23] & y[26];
  assign P[23][27] = x[23] & y[27];
  assign P[23][28] = x[23] & y[28];
  assign P[23][29] = x[23] & y[29];
  assign P[23][30] = x[23] & y[30];
  assign P[23][31] = x[23] & y[31];
  assign P[24][0] = x[24] & y[0];
  assign P[24][1] = x[24] & y[1];
  assign P[24][2] = x[24] & y[2];
  assign P[24][3] = x[24] & y[3];
  assign P[24][4] = x[24] & y[4];
  assign P[24][5] = x[24] & y[5];
  assign P[24][6] = x[24] & y[6];
  assign P[24][7] = x[24] & y[7];
  assign P[24][8] = x[24] & y[8];
  assign P[24][9] = x[24] & y[9];
  assign P[24][10] = x[24] & y[10];
  assign P[24][11] = x[24] & y[11];
  assign P[24][12] = x[24] & y[12];
  assign P[24][13] = x[24] & y[13];
  assign P[24][14] = x[24] & y[14];
  assign P[24][15] = x[24] & y[15];
  assign P[24][16] = x[24] & y[16];
  assign P[24][17] = x[24] & y[17];
  assign P[24][18] = x[24] & y[18];
  assign P[24][19] = x[24] & y[19];
  assign P[24][20] = x[24] & y[20];
  assign P[24][21] = x[24] & y[21];
  assign P[24][22] = x[24] & y[22];
  assign P[24][23] = x[24] & y[23];
  assign P[24][24] = x[24] & y[24];
  assign P[24][25] = x[24] & y[25];
  assign P[24][26] = x[24] & y[26];
  assign P[24][27] = x[24] & y[27];
  assign P[24][28] = x[24] & y[28];
  assign P[24][29] = x[24] & y[29];
  assign P[24][30] = x[24] & y[30];
  assign P[24][31] = x[24] & y[31];
  assign P[25][0] = x[25] & y[0];
  assign P[25][1] = x[25] & y[1];
  assign P[25][2] = x[25] & y[2];
  assign P[25][3] = x[25] & y[3];
  assign P[25][4] = x[25] & y[4];
  assign P[25][5] = x[25] & y[5];
  assign P[25][6] = x[25] & y[6];
  assign P[25][7] = x[25] & y[7];
  assign P[25][8] = x[25] & y[8];
  assign P[25][9] = x[25] & y[9];
  assign P[25][10] = x[25] & y[10];
  assign P[25][11] = x[25] & y[11];
  assign P[25][12] = x[25] & y[12];
  assign P[25][13] = x[25] & y[13];
  assign P[25][14] = x[25] & y[14];
  assign P[25][15] = x[25] & y[15];
  assign P[25][16] = x[25] & y[16];
  assign P[25][17] = x[25] & y[17];
  assign P[25][18] = x[25] & y[18];
  assign P[25][19] = x[25] & y[19];
  assign P[25][20] = x[25] & y[20];
  assign P[25][21] = x[25] & y[21];
  assign P[25][22] = x[25] & y[22];
  assign P[25][23] = x[25] & y[23];
  assign P[25][24] = x[25] & y[24];
  assign P[25][25] = x[25] & y[25];
  assign P[25][26] = x[25] & y[26];
  assign P[25][27] = x[25] & y[27];
  assign P[25][28] = x[25] & y[28];
  assign P[25][29] = x[25] & y[29];
  assign P[25][30] = x[25] & y[30];
  assign P[25][31] = x[25] & y[31];
  assign P[26][0] = x[26] & y[0];
  assign P[26][1] = x[26] & y[1];
  assign P[26][2] = x[26] & y[2];
  assign P[26][3] = x[26] & y[3];
  assign P[26][4] = x[26] & y[4];
  assign P[26][5] = x[26] & y[5];
  assign P[26][6] = x[26] & y[6];
  assign P[26][7] = x[26] & y[7];
  assign P[26][8] = x[26] & y[8];
  assign P[26][9] = x[26] & y[9];
  assign P[26][10] = x[26] & y[10];
  assign P[26][11] = x[26] & y[11];
  assign P[26][12] = x[26] & y[12];
  assign P[26][13] = x[26] & y[13];
  assign P[26][14] = x[26] & y[14];
  assign P[26][15] = x[26] & y[15];
  assign P[26][16] = x[26] & y[16];
  assign P[26][17] = x[26] & y[17];
  assign P[26][18] = x[26] & y[18];
  assign P[26][19] = x[26] & y[19];
  assign P[26][20] = x[26] & y[20];
  assign P[26][21] = x[26] & y[21];
  assign P[26][22] = x[26] & y[22];
  assign P[26][23] = x[26] & y[23];
  assign P[26][24] = x[26] & y[24];
  assign P[26][25] = x[26] & y[25];
  assign P[26][26] = x[26] & y[26];
  assign P[26][27] = x[26] & y[27];
  assign P[26][28] = x[26] & y[28];
  assign P[26][29] = x[26] & y[29];
  assign P[26][30] = x[26] & y[30];
  assign P[26][31] = x[26] & y[31];
  assign P[27][0] = x[27] & y[0];
  assign P[27][1] = x[27] & y[1];
  assign P[27][2] = x[27] & y[2];
  assign P[27][3] = x[27] & y[3];
  assign P[27][4] = x[27] & y[4];
  assign P[27][5] = x[27] & y[5];
  assign P[27][6] = x[27] & y[6];
  assign P[27][7] = x[27] & y[7];
  assign P[27][8] = x[27] & y[8];
  assign P[27][9] = x[27] & y[9];
  assign P[27][10] = x[27] & y[10];
  assign P[27][11] = x[27] & y[11];
  assign P[27][12] = x[27] & y[12];
  assign P[27][13] = x[27] & y[13];
  assign P[27][14] = x[27] & y[14];
  assign P[27][15] = x[27] & y[15];
  assign P[27][16] = x[27] & y[16];
  assign P[27][17] = x[27] & y[17];
  assign P[27][18] = x[27] & y[18];
  assign P[27][19] = x[27] & y[19];
  assign P[27][20] = x[27] & y[20];
  assign P[27][21] = x[27] & y[21];
  assign P[27][22] = x[27] & y[22];
  assign P[27][23] = x[27] & y[23];
  assign P[27][24] = x[27] & y[24];
  assign P[27][25] = x[27] & y[25];
  assign P[27][26] = x[27] & y[26];
  assign P[27][27] = x[27] & y[27];
  assign P[27][28] = x[27] & y[28];
  assign P[27][29] = x[27] & y[29];
  assign P[27][30] = x[27] & y[30];
  assign P[27][31] = x[27] & y[31];
  assign P[28][0] = x[28] & y[0];
  assign P[28][1] = x[28] & y[1];
  assign P[28][2] = x[28] & y[2];
  assign P[28][3] = x[28] & y[3];
  assign P[28][4] = x[28] & y[4];
  assign P[28][5] = x[28] & y[5];
  assign P[28][6] = x[28] & y[6];
  assign P[28][7] = x[28] & y[7];
  assign P[28][8] = x[28] & y[8];
  assign P[28][9] = x[28] & y[9];
  assign P[28][10] = x[28] & y[10];
  assign P[28][11] = x[28] & y[11];
  assign P[28][12] = x[28] & y[12];
  assign P[28][13] = x[28] & y[13];
  assign P[28][14] = x[28] & y[14];
  assign P[28][15] = x[28] & y[15];
  assign P[28][16] = x[28] & y[16];
  assign P[28][17] = x[28] & y[17];
  assign P[28][18] = x[28] & y[18];
  assign P[28][19] = x[28] & y[19];
  assign P[28][20] = x[28] & y[20];
  assign P[28][21] = x[28] & y[21];
  assign P[28][22] = x[28] & y[22];
  assign P[28][23] = x[28] & y[23];
  assign P[28][24] = x[28] & y[24];
  assign P[28][25] = x[28] & y[25];
  assign P[28][26] = x[28] & y[26];
  assign P[28][27] = x[28] & y[27];
  assign P[28][28] = x[28] & y[28];
  assign P[28][29] = x[28] & y[29];
  assign P[28][30] = x[28] & y[30];
  assign P[28][31] = x[28] & y[31];
  assign P[29][0] = x[29] & y[0];
  assign P[29][1] = x[29] & y[1];
  assign P[29][2] = x[29] & y[2];
  assign P[29][3] = x[29] & y[3];
  assign P[29][4] = x[29] & y[4];
  assign P[29][5] = x[29] & y[5];
  assign P[29][6] = x[29] & y[6];
  assign P[29][7] = x[29] & y[7];
  assign P[29][8] = x[29] & y[8];
  assign P[29][9] = x[29] & y[9];
  assign P[29][10] = x[29] & y[10];
  assign P[29][11] = x[29] & y[11];
  assign P[29][12] = x[29] & y[12];
  assign P[29][13] = x[29] & y[13];
  assign P[29][14] = x[29] & y[14];
  assign P[29][15] = x[29] & y[15];
  assign P[29][16] = x[29] & y[16];
  assign P[29][17] = x[29] & y[17];
  assign P[29][18] = x[29] & y[18];
  assign P[29][19] = x[29] & y[19];
  assign P[29][20] = x[29] & y[20];
  assign P[29][21] = x[29] & y[21];
  assign P[29][22] = x[29] & y[22];
  assign P[29][23] = x[29] & y[23];
  assign P[29][24] = x[29] & y[24];
  assign P[29][25] = x[29] & y[25];
  assign P[29][26] = x[29] & y[26];
  assign P[29][27] = x[29] & y[27];
  assign P[29][28] = x[29] & y[28];
  assign P[29][29] = x[29] & y[29];
  assign P[29][30] = x[29] & y[30];
  assign P[29][31] = x[29] & y[31];
  assign P[30][0] = x[30] & y[0];
  assign P[30][1] = x[30] & y[1];
  assign P[30][2] = x[30] & y[2];
  assign P[30][3] = x[30] & y[3];
  assign P[30][4] = x[30] & y[4];
  assign P[30][5] = x[30] & y[5];
  assign P[30][6] = x[30] & y[6];
  assign P[30][7] = x[30] & y[7];
  assign P[30][8] = x[30] & y[8];
  assign P[30][9] = x[30] & y[9];
  assign P[30][10] = x[30] & y[10];
  assign P[30][11] = x[30] & y[11];
  assign P[30][12] = x[30] & y[12];
  assign P[30][13] = x[30] & y[13];
  assign P[30][14] = x[30] & y[14];
  assign P[30][15] = x[30] & y[15];
  assign P[30][16] = x[30] & y[16];
  assign P[30][17] = x[30] & y[17];
  assign P[30][18] = x[30] & y[18];
  assign P[30][19] = x[30] & y[19];
  assign P[30][20] = x[30] & y[20];
  assign P[30][21] = x[30] & y[21];
  assign P[30][22] = x[30] & y[22];
  assign P[30][23] = x[30] & y[23];
  assign P[30][24] = x[30] & y[24];
  assign P[30][25] = x[30] & y[25];
  assign P[30][26] = x[30] & y[26];
  assign P[30][27] = x[30] & y[27];
  assign P[30][28] = x[30] & y[28];
  assign P[30][29] = x[30] & y[29];
  assign P[30][30] = x[30] & y[30];
  assign P[30][31] = x[30] & y[31];
  assign P[31][0] = x[31] & y[0];
  assign P[31][1] = x[31] & y[1];
  assign P[31][2] = x[31] & y[2];
  assign P[31][3] = x[31] & y[3];
  assign P[31][4] = x[31] & y[4];
  assign P[31][5] = x[31] & y[5];
  assign P[31][6] = x[31] & y[6];
  assign P[31][7] = x[31] & y[7];
  assign P[31][8] = x[31] & y[8];
  assign P[31][9] = x[31] & y[9];
  assign P[31][10] = x[31] & y[10];
  assign P[31][11] = x[31] & y[11];
  assign P[31][12] = x[31] & y[12];
  assign P[31][13] = x[31] & y[13];
  assign P[31][14] = x[31] & y[14];
  assign P[31][15] = x[31] & y[15];
  assign P[31][16] = x[31] & y[16];
  assign P[31][17] = x[31] & y[17];
  assign P[31][18] = x[31] & y[18];
  assign P[31][19] = x[31] & y[19];
  assign P[31][20] = x[31] & y[20];
  assign P[31][21] = x[31] & y[21];
  assign P[31][22] = x[31] & y[22];
  assign P[31][23] = x[31] & y[23];
  assign P[31][24] = x[31] & y[24];
  assign P[31][25] = x[31] & y[25];
  assign P[31][26] = x[31] & y[26];
  assign P[31][27] = x[31] & y[27];
  assign P[31][28] = x[31] & y[28];
  assign P[31][29] = x[31] & y[29];
  assign P[31][30] = x[31] & y[30];
  assign P[31][31] = x[31] & y[31];

  ha HA_00000000 (P[1][31],P[2][30],S[0],C[0]);
  fa FA_00000001 (P[0][31],P[1][30],P[2][29],S[1],C[1]);
  fa FA_00000002 (P[0][30],P[1][29],P[2][28],S[2],C[2]);
  fa FA_00000003 (P[0][29],P[1][28],P[2][27],S[3],C[3]);
  fa FA_00000004 (P[0][28],P[1][27],P[2][26],S[4],C[4]);
  fa FA_00000005 (P[0][27],P[1][26],P[2][25],S[5],C[5]);
  fa FA_00000006 (P[0][26],P[1][25],P[2][24],S[6],C[6]);
  fa FA_00000007 (P[0][25],P[1][24],P[2][23],S[7],C[7]);
  fa FA_00000008 (P[0][24],P[1][23],P[2][22],S[8],C[8]);
  fa FA_00000009 (P[0][23],P[1][22],P[2][21],S[9],C[9]);
  fa FA_00000010 (P[0][22],P[1][21],P[2][20],S[10],C[10]);
  fa FA_00000011 (P[0][21],P[1][20],P[2][19],S[11],C[11]);
  fa FA_00000012 (P[0][20],P[1][19],P[2][18],S[12],C[12]);
  fa FA_00000013 (P[0][19],P[1][18],P[2][17],S[13],C[13]);
  fa FA_00000014 (P[0][18],P[1][17],P[2][16],S[14],C[14]);
  fa FA_00000015 (P[0][17],P[1][16],P[2][15],S[15],C[15]);
  fa FA_00000016 (P[0][16],P[1][15],P[2][14],S[16],C[16]);
  fa FA_00000017 (P[0][15],P[1][14],P[2][13],S[17],C[17]);
  fa FA_00000018 (P[0][14],P[1][13],P[2][12],S[18],C[18]);
  fa FA_00000019 (P[0][13],P[1][12],P[2][11],S[19],C[19]);
  fa FA_00000020 (P[0][12],P[1][11],P[2][10],S[20],C[20]);
  fa FA_00000021 (P[0][11],P[1][10],P[2][9],S[21],C[21]);
  fa FA_00000022 (P[0][10],P[1][9],P[2][8],S[22],C[22]);
  fa FA_00000023 (P[0][9],P[1][8],P[2][7],S[23],C[23]);
  fa FA_00000024 (P[0][8],P[1][7],P[2][6],S[24],C[24]);
  fa FA_00000025 (P[0][7],P[1][6],P[2][5],S[25],C[25]);
  fa FA_00000026 (P[0][6],P[1][5],P[2][4],S[26],C[26]);
  fa FA_00000027 (P[0][5],P[1][4],P[2][3],S[27],C[27]);
  fa FA_00000028 (P[0][4],P[1][3],P[2][2],S[28],C[28]);
  fa FA_00000029 (P[0][3],P[1][2],P[2][1],S[29],C[29]);
  fa FA_00000030 (P[0][2],P[1][1],P[2][0],S[30],C[30]);
  ha HA_00000031 (P[0][1],P[1][0],S[31],C[31]);
  ha HA_00000032 (P[4][31],P[5][30],S[32],C[32]);
  fa FA_00000033 (P[3][31],P[4][30],P[5][29],S[33],C[33]);
  fa FA_00000034 (P[3][30],P[4][29],P[5][28],S[34],C[34]);
  fa FA_00000035 (P[3][29],P[4][28],P[5][27],S[35],C[35]);
  fa FA_00000036 (P[3][28],P[4][27],P[5][26],S[36],C[36]);
  fa FA_00000037 (P[3][27],P[4][26],P[5][25],S[37],C[37]);
  fa FA_00000038 (P[3][26],P[4][25],P[5][24],S[38],C[38]);
  fa FA_00000039 (P[3][25],P[4][24],P[5][23],S[39],C[39]);
  fa FA_00000040 (P[3][24],P[4][23],P[5][22],S[40],C[40]);
  fa FA_00000041 (P[3][23],P[4][22],P[5][21],S[41],C[41]);
  fa FA_00000042 (P[3][22],P[4][21],P[5][20],S[42],C[42]);
  fa FA_00000043 (P[3][21],P[4][20],P[5][19],S[43],C[43]);
  fa FA_00000044 (P[3][20],P[4][19],P[5][18],S[44],C[44]);
  fa FA_00000045 (P[3][19],P[4][18],P[5][17],S[45],C[45]);
  fa FA_00000046 (P[3][18],P[4][17],P[5][16],S[46],C[46]);
  fa FA_00000047 (P[3][17],P[4][16],P[5][15],S[47],C[47]);
  fa FA_00000048 (P[3][16],P[4][15],P[5][14],S[48],C[48]);
  fa FA_00000049 (P[3][15],P[4][14],P[5][13],S[49],C[49]);
  fa FA_00000050 (P[3][14],P[4][13],P[5][12],S[50],C[50]);
  fa FA_00000051 (P[3][13],P[4][12],P[5][11],S[51],C[51]);
  fa FA_00000052 (P[3][12],P[4][11],P[5][10],S[52],C[52]);
  fa FA_00000053 (P[3][11],P[4][10],P[5][9],S[53],C[53]);
  fa FA_00000054 (P[3][10],P[4][9],P[5][8],S[54],C[54]);
  fa FA_00000055 (P[3][9],P[4][8],P[5][7],S[55],C[55]);
  fa FA_00000056 (P[3][8],P[4][7],P[5][6],S[56],C[56]);
  fa FA_00000057 (P[3][7],P[4][6],P[5][5],S[57],C[57]);
  fa FA_00000058 (P[3][6],P[4][5],P[5][4],S[58],C[58]);
  fa FA_00000059 (P[3][5],P[4][4],P[5][3],S[59],C[59]);
  fa FA_00000060 (P[3][4],P[4][3],P[5][2],S[60],C[60]);
  fa FA_00000061 (P[3][3],P[4][2],P[5][1],S[61],C[61]);
  fa FA_00000062 (P[3][2],P[4][1],P[5][0],S[62],C[62]);
  ha HA_00000063 (P[3][1],P[4][0],S[63],C[63]);
  ha HA_00000064 (P[7][31],P[8][30],S[64],C[64]);
  fa FA_00000065 (P[6][31],P[7][30],P[8][29],S[65],C[65]);
  fa FA_00000066 (P[6][30],P[7][29],P[8][28],S[66],C[66]);
  fa FA_00000067 (P[6][29],P[7][28],P[8][27],S[67],C[67]);
  fa FA_00000068 (P[6][28],P[7][27],P[8][26],S[68],C[68]);
  fa FA_00000069 (P[6][27],P[7][26],P[8][25],S[69],C[69]);
  fa FA_00000070 (P[6][26],P[7][25],P[8][24],S[70],C[70]);
  fa FA_00000071 (P[6][25],P[7][24],P[8][23],S[71],C[71]);
  fa FA_00000072 (P[6][24],P[7][23],P[8][22],S[72],C[72]);
  fa FA_00000073 (P[6][23],P[7][22],P[8][21],S[73],C[73]);
  fa FA_00000074 (P[6][22],P[7][21],P[8][20],S[74],C[74]);
  fa FA_00000075 (P[6][21],P[7][20],P[8][19],S[75],C[75]);
  fa FA_00000076 (P[6][20],P[7][19],P[8][18],S[76],C[76]);
  fa FA_00000077 (P[6][19],P[7][18],P[8][17],S[77],C[77]);
  fa FA_00000078 (P[6][18],P[7][17],P[8][16],S[78],C[78]);
  fa FA_00000079 (P[6][17],P[7][16],P[8][15],S[79],C[79]);
  fa FA_00000080 (P[6][16],P[7][15],P[8][14],S[80],C[80]);
  fa FA_00000081 (P[6][15],P[7][14],P[8][13],S[81],C[81]);
  fa FA_00000082 (P[6][14],P[7][13],P[8][12],S[82],C[82]);
  fa FA_00000083 (P[6][13],P[7][12],P[8][11],S[83],C[83]);
  fa FA_00000084 (P[6][12],P[7][11],P[8][10],S[84],C[84]);
  fa FA_00000085 (P[6][11],P[7][10],P[8][9],S[85],C[85]);
  fa FA_00000086 (P[6][10],P[7][9],P[8][8],S[86],C[86]);
  fa FA_00000087 (P[6][9],P[7][8],P[8][7],S[87],C[87]);
  fa FA_00000088 (P[6][8],P[7][7],P[8][6],S[88],C[88]);
  fa FA_00000089 (P[6][7],P[7][6],P[8][5],S[89],C[89]);
  fa FA_00000090 (P[6][6],P[7][5],P[8][4],S[90],C[90]);
  fa FA_00000091 (P[6][5],P[7][4],P[8][3],S[91],C[91]);
  fa FA_00000092 (P[6][4],P[7][3],P[8][2],S[92],C[92]);
  fa FA_00000093 (P[6][3],P[7][2],P[8][1],S[93],C[93]);
  fa FA_00000094 (P[6][2],P[7][1],P[8][0],S[94],C[94]);
  ha HA_00000095 (P[6][1],P[7][0],S[95],C[95]);
  ha HA_00000096 (P[10][31],P[11][30],S[96],C[96]);
  fa FA_00000097 (P[9][31],P[10][30],P[11][29],S[97],C[97]);
  fa FA_00000098 (P[9][30],P[10][29],P[11][28],S[98],C[98]);
  fa FA_00000099 (P[9][29],P[10][28],P[11][27],S[99],C[99]);
  fa FA_00000100 (P[9][28],P[10][27],P[11][26],S[100],C[100]);
  fa FA_00000101 (P[9][27],P[10][26],P[11][25],S[101],C[101]);
  fa FA_00000102 (P[9][26],P[10][25],P[11][24],S[102],C[102]);
  fa FA_00000103 (P[9][25],P[10][24],P[11][23],S[103],C[103]);
  fa FA_00000104 (P[9][24],P[10][23],P[11][22],S[104],C[104]);
  fa FA_00000105 (P[9][23],P[10][22],P[11][21],S[105],C[105]);
  fa FA_00000106 (P[9][22],P[10][21],P[11][20],S[106],C[106]);
  fa FA_00000107 (P[9][21],P[10][20],P[11][19],S[107],C[107]);
  fa FA_00000108 (P[9][20],P[10][19],P[11][18],S[108],C[108]);
  fa FA_00000109 (P[9][19],P[10][18],P[11][17],S[109],C[109]);
  fa FA_00000110 (P[9][18],P[10][17],P[11][16],S[110],C[110]);
  fa FA_00000111 (P[9][17],P[10][16],P[11][15],S[111],C[111]);
  fa FA_00000112 (P[9][16],P[10][15],P[11][14],S[112],C[112]);
  fa FA_00000113 (P[9][15],P[10][14],P[11][13],S[113],C[113]);
  fa FA_00000114 (P[9][14],P[10][13],P[11][12],S[114],C[114]);
  fa FA_00000115 (P[9][13],P[10][12],P[11][11],S[115],C[115]);
  fa FA_00000116 (P[9][12],P[10][11],P[11][10],S[116],C[116]);
  fa FA_00000117 (P[9][11],P[10][10],P[11][9],S[117],C[117]);
  fa FA_00000118 (P[9][10],P[10][9],P[11][8],S[118],C[118]);
  fa FA_00000119 (P[9][9],P[10][8],P[11][7],S[119],C[119]);
  fa FA_00000120 (P[9][8],P[10][7],P[11][6],S[120],C[120]);
  fa FA_00000121 (P[9][7],P[10][6],P[11][5],S[121],C[121]);
  fa FA_00000122 (P[9][6],P[10][5],P[11][4],S[122],C[122]);
  fa FA_00000123 (P[9][5],P[10][4],P[11][3],S[123],C[123]);
  fa FA_00000124 (P[9][4],P[10][3],P[11][2],S[124],C[124]);
  fa FA_00000125 (P[9][3],P[10][2],P[11][1],S[125],C[125]);
  fa FA_00000126 (P[9][2],P[10][1],P[11][0],S[126],C[126]);
  ha HA_00000127 (P[9][1],P[10][0],S[127],C[127]);
  ha HA_00000128 (P[13][31],P[14][30],S[128],C[128]);
  fa FA_00000129 (P[12][31],P[13][30],P[14][29],S[129],C[129]);
  fa FA_00000130 (P[12][30],P[13][29],P[14][28],S[130],C[130]);
  fa FA_00000131 (P[12][29],P[13][28],P[14][27],S[131],C[131]);
  fa FA_00000132 (P[12][28],P[13][27],P[14][26],S[132],C[132]);
  fa FA_00000133 (P[12][27],P[13][26],P[14][25],S[133],C[133]);
  fa FA_00000134 (P[12][26],P[13][25],P[14][24],S[134],C[134]);
  fa FA_00000135 (P[12][25],P[13][24],P[14][23],S[135],C[135]);
  fa FA_00000136 (P[12][24],P[13][23],P[14][22],S[136],C[136]);
  fa FA_00000137 (P[12][23],P[13][22],P[14][21],S[137],C[137]);
  fa FA_00000138 (P[12][22],P[13][21],P[14][20],S[138],C[138]);
  fa FA_00000139 (P[12][21],P[13][20],P[14][19],S[139],C[139]);
  fa FA_00000140 (P[12][20],P[13][19],P[14][18],S[140],C[140]);
  fa FA_00000141 (P[12][19],P[13][18],P[14][17],S[141],C[141]);
  fa FA_00000142 (P[12][18],P[13][17],P[14][16],S[142],C[142]);
  fa FA_00000143 (P[12][17],P[13][16],P[14][15],S[143],C[143]);
  fa FA_00000144 (P[12][16],P[13][15],P[14][14],S[144],C[144]);
  fa FA_00000145 (P[12][15],P[13][14],P[14][13],S[145],C[145]);
  fa FA_00000146 (P[12][14],P[13][13],P[14][12],S[146],C[146]);
  fa FA_00000147 (P[12][13],P[13][12],P[14][11],S[147],C[147]);
  fa FA_00000148 (P[12][12],P[13][11],P[14][10],S[148],C[148]);
  fa FA_00000149 (P[12][11],P[13][10],P[14][9],S[149],C[149]);
  fa FA_00000150 (P[12][10],P[13][9],P[14][8],S[150],C[150]);
  fa FA_00000151 (P[12][9],P[13][8],P[14][7],S[151],C[151]);
  fa FA_00000152 (P[12][8],P[13][7],P[14][6],S[152],C[152]);
  fa FA_00000153 (P[12][7],P[13][6],P[14][5],S[153],C[153]);
  fa FA_00000154 (P[12][6],P[13][5],P[14][4],S[154],C[154]);
  fa FA_00000155 (P[12][5],P[13][4],P[14][3],S[155],C[155]);
  fa FA_00000156 (P[12][4],P[13][3],P[14][2],S[156],C[156]);
  fa FA_00000157 (P[12][3],P[13][2],P[14][1],S[157],C[157]);
  fa FA_00000158 (P[12][2],P[13][1],P[14][0],S[158],C[158]);
  ha HA_00000159 (P[12][1],P[13][0],S[159],C[159]);
  ha HA_00000160 (P[16][31],P[17][30],S[160],C[160]);
  fa FA_00000161 (P[15][31],P[16][30],P[17][29],S[161],C[161]);
  fa FA_00000162 (P[15][30],P[16][29],P[17][28],S[162],C[162]);
  fa FA_00000163 (P[15][29],P[16][28],P[17][27],S[163],C[163]);
  fa FA_00000164 (P[15][28],P[16][27],P[17][26],S[164],C[164]);
  fa FA_00000165 (P[15][27],P[16][26],P[17][25],S[165],C[165]);
  fa FA_00000166 (P[15][26],P[16][25],P[17][24],S[166],C[166]);
  fa FA_00000167 (P[15][25],P[16][24],P[17][23],S[167],C[167]);
  fa FA_00000168 (P[15][24],P[16][23],P[17][22],S[168],C[168]);
  fa FA_00000169 (P[15][23],P[16][22],P[17][21],S[169],C[169]);
  fa FA_00000170 (P[15][22],P[16][21],P[17][20],S[170],C[170]);
  fa FA_00000171 (P[15][21],P[16][20],P[17][19],S[171],C[171]);
  fa FA_00000172 (P[15][20],P[16][19],P[17][18],S[172],C[172]);
  fa FA_00000173 (P[15][19],P[16][18],P[17][17],S[173],C[173]);
  fa FA_00000174 (P[15][18],P[16][17],P[17][16],S[174],C[174]);
  fa FA_00000175 (P[15][17],P[16][16],P[17][15],S[175],C[175]);
  fa FA_00000176 (P[15][16],P[16][15],P[17][14],S[176],C[176]);
  fa FA_00000177 (P[15][15],P[16][14],P[17][13],S[177],C[177]);
  fa FA_00000178 (P[15][14],P[16][13],P[17][12],S[178],C[178]);
  fa FA_00000179 (P[15][13],P[16][12],P[17][11],S[179],C[179]);
  fa FA_00000180 (P[15][12],P[16][11],P[17][10],S[180],C[180]);
  fa FA_00000181 (P[15][11],P[16][10],P[17][9],S[181],C[181]);
  fa FA_00000182 (P[15][10],P[16][9],P[17][8],S[182],C[182]);
  fa FA_00000183 (P[15][9],P[16][8],P[17][7],S[183],C[183]);
  fa FA_00000184 (P[15][8],P[16][7],P[17][6],S[184],C[184]);
  fa FA_00000185 (P[15][7],P[16][6],P[17][5],S[185],C[185]);
  fa FA_00000186 (P[15][6],P[16][5],P[17][4],S[186],C[186]);
  fa FA_00000187 (P[15][5],P[16][4],P[17][3],S[187],C[187]);
  fa FA_00000188 (P[15][4],P[16][3],P[17][2],S[188],C[188]);
  fa FA_00000189 (P[15][3],P[16][2],P[17][1],S[189],C[189]);
  fa FA_00000190 (P[15][2],P[16][1],P[17][0],S[190],C[190]);
  ha HA_00000191 (P[15][1],P[16][0],S[191],C[191]);
  ha HA_00000192 (P[19][31],P[20][30],S[192],C[192]);
  fa FA_00000193 (P[18][31],P[19][30],P[20][29],S[193],C[193]);
  fa FA_00000194 (P[18][30],P[19][29],P[20][28],S[194],C[194]);
  fa FA_00000195 (P[18][29],P[19][28],P[20][27],S[195],C[195]);
  fa FA_00000196 (P[18][28],P[19][27],P[20][26],S[196],C[196]);
  fa FA_00000197 (P[18][27],P[19][26],P[20][25],S[197],C[197]);
  fa FA_00000198 (P[18][26],P[19][25],P[20][24],S[198],C[198]);
  fa FA_00000199 (P[18][25],P[19][24],P[20][23],S[199],C[199]);
  fa FA_00000200 (P[18][24],P[19][23],P[20][22],S[200],C[200]);
  fa FA_00000201 (P[18][23],P[19][22],P[20][21],S[201],C[201]);
  fa FA_00000202 (P[18][22],P[19][21],P[20][20],S[202],C[202]);
  fa FA_00000203 (P[18][21],P[19][20],P[20][19],S[203],C[203]);
  fa FA_00000204 (P[18][20],P[19][19],P[20][18],S[204],C[204]);
  fa FA_00000205 (P[18][19],P[19][18],P[20][17],S[205],C[205]);
  fa FA_00000206 (P[18][18],P[19][17],P[20][16],S[206],C[206]);
  fa FA_00000207 (P[18][17],P[19][16],P[20][15],S[207],C[207]);
  fa FA_00000208 (P[18][16],P[19][15],P[20][14],S[208],C[208]);
  fa FA_00000209 (P[18][15],P[19][14],P[20][13],S[209],C[209]);
  fa FA_00000210 (P[18][14],P[19][13],P[20][12],S[210],C[210]);
  fa FA_00000211 (P[18][13],P[19][12],P[20][11],S[211],C[211]);
  fa FA_00000212 (P[18][12],P[19][11],P[20][10],S[212],C[212]);
  fa FA_00000213 (P[18][11],P[19][10],P[20][9],S[213],C[213]);
  fa FA_00000214 (P[18][10],P[19][9],P[20][8],S[214],C[214]);
  fa FA_00000215 (P[18][9],P[19][8],P[20][7],S[215],C[215]);
  fa FA_00000216 (P[18][8],P[19][7],P[20][6],S[216],C[216]);
  fa FA_00000217 (P[18][7],P[19][6],P[20][5],S[217],C[217]);
  fa FA_00000218 (P[18][6],P[19][5],P[20][4],S[218],C[218]);
  fa FA_00000219 (P[18][5],P[19][4],P[20][3],S[219],C[219]);
  fa FA_00000220 (P[18][4],P[19][3],P[20][2],S[220],C[220]);
  fa FA_00000221 (P[18][3],P[19][2],P[20][1],S[221],C[221]);
  fa FA_00000222 (P[18][2],P[19][1],P[20][0],S[222],C[222]);
  ha HA_00000223 (P[18][1],P[19][0],S[223],C[223]);
  ha HA_00000224 (P[22][31],P[23][30],S[224],C[224]);
  fa FA_00000225 (P[21][31],P[22][30],P[23][29],S[225],C[225]);
  fa FA_00000226 (P[21][30],P[22][29],P[23][28],S[226],C[226]);
  fa FA_00000227 (P[21][29],P[22][28],P[23][27],S[227],C[227]);
  fa FA_00000228 (P[21][28],P[22][27],P[23][26],S[228],C[228]);
  fa FA_00000229 (P[21][27],P[22][26],P[23][25],S[229],C[229]);
  fa FA_00000230 (P[21][26],P[22][25],P[23][24],S[230],C[230]);
  fa FA_00000231 (P[21][25],P[22][24],P[23][23],S[231],C[231]);
  fa FA_00000232 (P[21][24],P[22][23],P[23][22],S[232],C[232]);
  fa FA_00000233 (P[21][23],P[22][22],P[23][21],S[233],C[233]);
  fa FA_00000234 (P[21][22],P[22][21],P[23][20],S[234],C[234]);
  fa FA_00000235 (P[21][21],P[22][20],P[23][19],S[235],C[235]);
  fa FA_00000236 (P[21][20],P[22][19],P[23][18],S[236],C[236]);
  fa FA_00000237 (P[21][19],P[22][18],P[23][17],S[237],C[237]);
  fa FA_00000238 (P[21][18],P[22][17],P[23][16],S[238],C[238]);
  fa FA_00000239 (P[21][17],P[22][16],P[23][15],S[239],C[239]);
  fa FA_00000240 (P[21][16],P[22][15],P[23][14],S[240],C[240]);
  fa FA_00000241 (P[21][15],P[22][14],P[23][13],S[241],C[241]);
  fa FA_00000242 (P[21][14],P[22][13],P[23][12],S[242],C[242]);
  fa FA_00000243 (P[21][13],P[22][12],P[23][11],S[243],C[243]);
  fa FA_00000244 (P[21][12],P[22][11],P[23][10],S[244],C[244]);
  fa FA_00000245 (P[21][11],P[22][10],P[23][9],S[245],C[245]);
  fa FA_00000246 (P[21][10],P[22][9],P[23][8],S[246],C[246]);
  fa FA_00000247 (P[21][9],P[22][8],P[23][7],S[247],C[247]);
  fa FA_00000248 (P[21][8],P[22][7],P[23][6],S[248],C[248]);
  fa FA_00000249 (P[21][7],P[22][6],P[23][5],S[249],C[249]);
  fa FA_00000250 (P[21][6],P[22][5],P[23][4],S[250],C[250]);
  fa FA_00000251 (P[21][5],P[22][4],P[23][3],S[251],C[251]);
  fa FA_00000252 (P[21][4],P[22][3],P[23][2],S[252],C[252]);
  fa FA_00000253 (P[21][3],P[22][2],P[23][1],S[253],C[253]);
  fa FA_00000254 (P[21][2],P[22][1],P[23][0],S[254],C[254]);
  ha HA_00000255 (P[21][1],P[22][0],S[255],C[255]);
  ha HA_00000256 (P[25][31],P[26][30],S[256],C[256]);
  fa FA_00000257 (P[24][31],P[25][30],P[26][29],S[257],C[257]);
  fa FA_00000258 (P[24][30],P[25][29],P[26][28],S[258],C[258]);
  fa FA_00000259 (P[24][29],P[25][28],P[26][27],S[259],C[259]);
  fa FA_00000260 (P[24][28],P[25][27],P[26][26],S[260],C[260]);
  fa FA_00000261 (P[24][27],P[25][26],P[26][25],S[261],C[261]);
  fa FA_00000262 (P[24][26],P[25][25],P[26][24],S[262],C[262]);
  fa FA_00000263 (P[24][25],P[25][24],P[26][23],S[263],C[263]);
  fa FA_00000264 (P[24][24],P[25][23],P[26][22],S[264],C[264]);
  fa FA_00000265 (P[24][23],P[25][22],P[26][21],S[265],C[265]);
  fa FA_00000266 (P[24][22],P[25][21],P[26][20],S[266],C[266]);
  fa FA_00000267 (P[24][21],P[25][20],P[26][19],S[267],C[267]);
  fa FA_00000268 (P[24][20],P[25][19],P[26][18],S[268],C[268]);
  fa FA_00000269 (P[24][19],P[25][18],P[26][17],S[269],C[269]);
  fa FA_00000270 (P[24][18],P[25][17],P[26][16],S[270],C[270]);
  fa FA_00000271 (P[24][17],P[25][16],P[26][15],S[271],C[271]);
  fa FA_00000272 (P[24][16],P[25][15],P[26][14],S[272],C[272]);
  fa FA_00000273 (P[24][15],P[25][14],P[26][13],S[273],C[273]);
  fa FA_00000274 (P[24][14],P[25][13],P[26][12],S[274],C[274]);
  fa FA_00000275 (P[24][13],P[25][12],P[26][11],S[275],C[275]);
  fa FA_00000276 (P[24][12],P[25][11],P[26][10],S[276],C[276]);
  fa FA_00000277 (P[24][11],P[25][10],P[26][9],S[277],C[277]);
  fa FA_00000278 (P[24][10],P[25][9],P[26][8],S[278],C[278]);
  fa FA_00000279 (P[24][9],P[25][8],P[26][7],S[279],C[279]);
  fa FA_00000280 (P[24][8],P[25][7],P[26][6],S[280],C[280]);
  fa FA_00000281 (P[24][7],P[25][6],P[26][5],S[281],C[281]);
  fa FA_00000282 (P[24][6],P[25][5],P[26][4],S[282],C[282]);
  fa FA_00000283 (P[24][5],P[25][4],P[26][3],S[283],C[283]);
  fa FA_00000284 (P[24][4],P[25][3],P[26][2],S[284],C[284]);
  fa FA_00000285 (P[24][3],P[25][2],P[26][1],S[285],C[285]);
  fa FA_00000286 (P[24][2],P[25][1],P[26][0],S[286],C[286]);
  ha HA_00000287 (P[24][1],P[25][0],S[287],C[287]);
  ha HA_00000288 (P[28][31],P[29][30],S[288],C[288]);
  fa FA_00000289 (P[27][31],P[28][30],P[29][29],S[289],C[289]);
  fa FA_00000290 (P[27][30],P[28][29],P[29][28],S[290],C[290]);
  fa FA_00000291 (P[27][29],P[28][28],P[29][27],S[291],C[291]);
  fa FA_00000292 (P[27][28],P[28][27],P[29][26],S[292],C[292]);
  fa FA_00000293 (P[27][27],P[28][26],P[29][25],S[293],C[293]);
  fa FA_00000294 (P[27][26],P[28][25],P[29][24],S[294],C[294]);
  fa FA_00000295 (P[27][25],P[28][24],P[29][23],S[295],C[295]);
  fa FA_00000296 (P[27][24],P[28][23],P[29][22],S[296],C[296]);
  fa FA_00000297 (P[27][23],P[28][22],P[29][21],S[297],C[297]);
  fa FA_00000298 (P[27][22],P[28][21],P[29][20],S[298],C[298]);
  fa FA_00000299 (P[27][21],P[28][20],P[29][19],S[299],C[299]);
  fa FA_00000300 (P[27][20],P[28][19],P[29][18],S[300],C[300]);
  fa FA_00000301 (P[27][19],P[28][18],P[29][17],S[301],C[301]);
  fa FA_00000302 (P[27][18],P[28][17],P[29][16],S[302],C[302]);
  fa FA_00000303 (P[27][17],P[28][16],P[29][15],S[303],C[303]);
  fa FA_00000304 (P[27][16],P[28][15],P[29][14],S[304],C[304]);
  fa FA_00000305 (P[27][15],P[28][14],P[29][13],S[305],C[305]);
  fa FA_00000306 (P[27][14],P[28][13],P[29][12],S[306],C[306]);
  fa FA_00000307 (P[27][13],P[28][12],P[29][11],S[307],C[307]);
  fa FA_00000308 (P[27][12],P[28][11],P[29][10],S[308],C[308]);
  fa FA_00000309 (P[27][11],P[28][10],P[29][9],S[309],C[309]);
  fa FA_00000310 (P[27][10],P[28][9],P[29][8],S[310],C[310]);
  fa FA_00000311 (P[27][9],P[28][8],P[29][7],S[311],C[311]);
  fa FA_00000312 (P[27][8],P[28][7],P[29][6],S[312],C[312]);
  fa FA_00000313 (P[27][7],P[28][6],P[29][5],S[313],C[313]);
  fa FA_00000314 (P[27][6],P[28][5],P[29][4],S[314],C[314]);
  fa FA_00000315 (P[27][5],P[28][4],P[29][3],S[315],C[315]);
  fa FA_00000316 (P[27][4],P[28][3],P[29][2],S[316],C[316]);
  fa FA_00000317 (P[27][3],P[28][2],P[29][1],S[317],C[317]);
  fa FA_00000318 (P[27][2],P[28][1],P[29][0],S[318],C[318]);
  ha HA_00000319 (P[27][1],P[28][0],S[319],C[319]);
  fa FA_00000320 (P[2][31],C[0],S[34],S[320],C[320]);
  fa FA_00000321 (S[0],C[1],S[35],S[321],C[321]);
  fa FA_00000322 (S[1],C[2],S[36],S[322],C[322]);
  fa FA_00000323 (S[2],C[3],S[37],S[323],C[323]);
  fa FA_00000324 (S[3],C[4],S[38],S[324],C[324]);
  fa FA_00000325 (S[4],C[5],S[39],S[325],C[325]);
  fa FA_00000326 (S[5],C[6],S[40],S[326],C[326]);
  fa FA_00000327 (S[6],C[7],S[41],S[327],C[327]);
  fa FA_00000328 (S[7],C[8],S[42],S[328],C[328]);
  fa FA_00000329 (S[8],C[9],S[43],S[329],C[329]);
  fa FA_00000330 (S[9],C[10],S[44],S[330],C[330]);
  fa FA_00000331 (S[10],C[11],S[45],S[331],C[331]);
  fa FA_00000332 (S[11],C[12],S[46],S[332],C[332]);
  fa FA_00000333 (S[12],C[13],S[47],S[333],C[333]);
  fa FA_00000334 (S[13],C[14],S[48],S[334],C[334]);
  fa FA_00000335 (S[14],C[15],S[49],S[335],C[335]);
  fa FA_00000336 (S[15],C[16],S[50],S[336],C[336]);
  fa FA_00000337 (S[16],C[17],S[51],S[337],C[337]);
  fa FA_00000338 (S[17],C[18],S[52],S[338],C[338]);
  fa FA_00000339 (S[18],C[19],S[53],S[339],C[339]);
  fa FA_00000340 (S[19],C[20],S[54],S[340],C[340]);
  fa FA_00000341 (S[20],C[21],S[55],S[341],C[341]);
  fa FA_00000342 (S[21],C[22],S[56],S[342],C[342]);
  fa FA_00000343 (S[22],C[23],S[57],S[343],C[343]);
  fa FA_00000344 (S[23],C[24],S[58],S[344],C[344]);
  fa FA_00000345 (S[24],C[25],S[59],S[345],C[345]);
  fa FA_00000346 (S[25],C[26],S[60],S[346],C[346]);
  fa FA_00000347 (S[26],C[27],S[61],S[347],C[347]);
  fa FA_00000348 (S[27],C[28],S[62],S[348],C[348]);
  fa FA_00000349 (S[28],C[29],S[63],S[349],C[349]);
  fa FA_00000350 (S[29],C[30],P[3][0],S[350],C[350]);
  ha HA_00000351 (S[30],C[31],S[351],C[351]);
  ha HA_00000352 (P[8][31],C[64],S[352],C[352]);
  ha HA_00000353 (S[64],C[65],S[353],C[353]);
  ha HA_00000354 (S[65],C[66],S[354],C[354]);
  fa FA_00000355 (C[32],S[66],C[67],S[355],C[355]);
  fa FA_00000356 (C[33],S[67],C[68],S[356],C[356]);
  fa FA_00000357 (C[34],S[68],C[69],S[357],C[357]);
  fa FA_00000358 (C[35],S[69],C[70],S[358],C[358]);
  fa FA_00000359 (C[36],S[70],C[71],S[359],C[359]);
  fa FA_00000360 (C[37],S[71],C[72],S[360],C[360]);
  fa FA_00000361 (C[38],S[72],C[73],S[361],C[361]);
  fa FA_00000362 (C[39],S[73],C[74],S[362],C[362]);
  fa FA_00000363 (C[40],S[74],C[75],S[363],C[363]);
  fa FA_00000364 (C[41],S[75],C[76],S[364],C[364]);
  fa FA_00000365 (C[42],S[76],C[77],S[365],C[365]);
  fa FA_00000366 (C[43],S[77],C[78],S[366],C[366]);
  fa FA_00000367 (C[44],S[78],C[79],S[367],C[367]);
  fa FA_00000368 (C[45],S[79],C[80],S[368],C[368]);
  fa FA_00000369 (C[46],S[80],C[81],S[369],C[369]);
  fa FA_00000370 (C[47],S[81],C[82],S[370],C[370]);
  fa FA_00000371 (C[48],S[82],C[83],S[371],C[371]);
  fa FA_00000372 (C[49],S[83],C[84],S[372],C[372]);
  fa FA_00000373 (C[50],S[84],C[85],S[373],C[373]);
  fa FA_00000374 (C[51],S[85],C[86],S[374],C[374]);
  fa FA_00000375 (C[52],S[86],C[87],S[375],C[375]);
  fa FA_00000376 (C[53],S[87],C[88],S[376],C[376]);
  fa FA_00000377 (C[54],S[88],C[89],S[377],C[377]);
  fa FA_00000378 (C[55],S[89],C[90],S[378],C[378]);
  fa FA_00000379 (C[56],S[90],C[91],S[379],C[379]);
  fa FA_00000380 (C[57],S[91],C[92],S[380],C[380]);
  fa FA_00000381 (C[58],S[92],C[93],S[381],C[381]);
  fa FA_00000382 (C[59],S[93],C[94],S[382],C[382]);
  fa FA_00000383 (C[60],S[94],C[95],S[383],C[383]);
  ha HA_00000384 (C[61],S[95],S[384],C[384]);
  ha HA_00000385 (C[62],P[6][0],S[385],C[385]);
  fa FA_00000386 (P[11][31],C[96],S[130],S[386],C[386]);
  fa FA_00000387 (S[96],C[97],S[131],S[387],C[387]);
  fa FA_00000388 (S[97],C[98],S[132],S[388],C[388]);
  fa FA_00000389 (S[98],C[99],S[133],S[389],C[389]);
  fa FA_00000390 (S[99],C[100],S[134],S[390],C[390]);
  fa FA_00000391 (S[100],C[101],S[135],S[391],C[391]);
  fa FA_00000392 (S[101],C[102],S[136],S[392],C[392]);
  fa FA_00000393 (S[102],C[103],S[137],S[393],C[393]);
  fa FA_00000394 (S[103],C[104],S[138],S[394],C[394]);
  fa FA_00000395 (S[104],C[105],S[139],S[395],C[395]);
  fa FA_00000396 (S[105],C[106],S[140],S[396],C[396]);
  fa FA_00000397 (S[106],C[107],S[141],S[397],C[397]);
  fa FA_00000398 (S[107],C[108],S[142],S[398],C[398]);
  fa FA_00000399 (S[108],C[109],S[143],S[399],C[399]);
  fa FA_00000400 (S[109],C[110],S[144],S[400],C[400]);
  fa FA_00000401 (S[110],C[111],S[145],S[401],C[401]);
  fa FA_00000402 (S[111],C[112],S[146],S[402],C[402]);
  fa FA_00000403 (S[112],C[113],S[147],S[403],C[403]);
  fa FA_00000404 (S[113],C[114],S[148],S[404],C[404]);
  fa FA_00000405 (S[114],C[115],S[149],S[405],C[405]);
  fa FA_00000406 (S[115],C[116],S[150],S[406],C[406]);
  fa FA_00000407 (S[116],C[117],S[151],S[407],C[407]);
  fa FA_00000408 (S[117],C[118],S[152],S[408],C[408]);
  fa FA_00000409 (S[118],C[119],S[153],S[409],C[409]);
  fa FA_00000410 (S[119],C[120],S[154],S[410],C[410]);
  fa FA_00000411 (S[120],C[121],S[155],S[411],C[411]);
  fa FA_00000412 (S[121],C[122],S[156],S[412],C[412]);
  fa FA_00000413 (S[122],C[123],S[157],S[413],C[413]);
  fa FA_00000414 (S[123],C[124],S[158],S[414],C[414]);
  fa FA_00000415 (S[124],C[125],S[159],S[415],C[415]);
  fa FA_00000416 (S[125],C[126],P[12][0],S[416],C[416]);
  ha HA_00000417 (S[126],C[127],S[417],C[417]);
  ha HA_00000418 (P[17][31],C[160],S[418],C[418]);
  ha HA_00000419 (S[160],C[161],S[419],C[419]);
  ha HA_00000420 (S[161],C[162],S[420],C[420]);
  fa FA_00000421 (C[128],S[162],C[163],S[421],C[421]);
  fa FA_00000422 (C[129],S[163],C[164],S[422],C[422]);
  fa FA_00000423 (C[130],S[164],C[165],S[423],C[423]);
  fa FA_00000424 (C[131],S[165],C[166],S[424],C[424]);
  fa FA_00000425 (C[132],S[166],C[167],S[425],C[425]);
  fa FA_00000426 (C[133],S[167],C[168],S[426],C[426]);
  fa FA_00000427 (C[134],S[168],C[169],S[427],C[427]);
  fa FA_00000428 (C[135],S[169],C[170],S[428],C[428]);
  fa FA_00000429 (C[136],S[170],C[171],S[429],C[429]);
  fa FA_00000430 (C[137],S[171],C[172],S[430],C[430]);
  fa FA_00000431 (C[138],S[172],C[173],S[431],C[431]);
  fa FA_00000432 (C[139],S[173],C[174],S[432],C[432]);
  fa FA_00000433 (C[140],S[174],C[175],S[433],C[433]);
  fa FA_00000434 (C[141],S[175],C[176],S[434],C[434]);
  fa FA_00000435 (C[142],S[176],C[177],S[435],C[435]);
  fa FA_00000436 (C[143],S[177],C[178],S[436],C[436]);
  fa FA_00000437 (C[144],S[178],C[179],S[437],C[437]);
  fa FA_00000438 (C[145],S[179],C[180],S[438],C[438]);
  fa FA_00000439 (C[146],S[180],C[181],S[439],C[439]);
  fa FA_00000440 (C[147],S[181],C[182],S[440],C[440]);
  fa FA_00000441 (C[148],S[182],C[183],S[441],C[441]);
  fa FA_00000442 (C[149],S[183],C[184],S[442],C[442]);
  fa FA_00000443 (C[150],S[184],C[185],S[443],C[443]);
  fa FA_00000444 (C[151],S[185],C[186],S[444],C[444]);
  fa FA_00000445 (C[152],S[186],C[187],S[445],C[445]);
  fa FA_00000446 (C[153],S[187],C[188],S[446],C[446]);
  fa FA_00000447 (C[154],S[188],C[189],S[447],C[447]);
  fa FA_00000448 (C[155],S[189],C[190],S[448],C[448]);
  fa FA_00000449 (C[156],S[190],C[191],S[449],C[449]);
  ha HA_00000450 (C[157],S[191],S[450],C[450]);
  ha HA_00000451 (C[158],P[15][0],S[451],C[451]);
  fa FA_00000452 (P[20][31],C[192],S[226],S[452],C[452]);
  fa FA_00000453 (S[192],C[193],S[227],S[453],C[453]);
  fa FA_00000454 (S[193],C[194],S[228],S[454],C[454]);
  fa FA_00000455 (S[194],C[195],S[229],S[455],C[455]);
  fa FA_00000456 (S[195],C[196],S[230],S[456],C[456]);
  fa FA_00000457 (S[196],C[197],S[231],S[457],C[457]);
  fa FA_00000458 (S[197],C[198],S[232],S[458],C[458]);
  fa FA_00000459 (S[198],C[199],S[233],S[459],C[459]);
  fa FA_00000460 (S[199],C[200],S[234],S[460],C[460]);
  fa FA_00000461 (S[200],C[201],S[235],S[461],C[461]);
  fa FA_00000462 (S[201],C[202],S[236],S[462],C[462]);
  fa FA_00000463 (S[202],C[203],S[237],S[463],C[463]);
  fa FA_00000464 (S[203],C[204],S[238],S[464],C[464]);
  fa FA_00000465 (S[204],C[205],S[239],S[465],C[465]);
  fa FA_00000466 (S[205],C[206],S[240],S[466],C[466]);
  fa FA_00000467 (S[206],C[207],S[241],S[467],C[467]);
  fa FA_00000468 (S[207],C[208],S[242],S[468],C[468]);
  fa FA_00000469 (S[208],C[209],S[243],S[469],C[469]);
  fa FA_00000470 (S[209],C[210],S[244],S[470],C[470]);
  fa FA_00000471 (S[210],C[211],S[245],S[471],C[471]);
  fa FA_00000472 (S[211],C[212],S[246],S[472],C[472]);
  fa FA_00000473 (S[212],C[213],S[247],S[473],C[473]);
  fa FA_00000474 (S[213],C[214],S[248],S[474],C[474]);
  fa FA_00000475 (S[214],C[215],S[249],S[475],C[475]);
  fa FA_00000476 (S[215],C[216],S[250],S[476],C[476]);
  fa FA_00000477 (S[216],C[217],S[251],S[477],C[477]);
  fa FA_00000478 (S[217],C[218],S[252],S[478],C[478]);
  fa FA_00000479 (S[218],C[219],S[253],S[479],C[479]);
  fa FA_00000480 (S[219],C[220],S[254],S[480],C[480]);
  fa FA_00000481 (S[220],C[221],S[255],S[481],C[481]);
  fa FA_00000482 (S[221],C[222],P[21][0],S[482],C[482]);
  ha HA_00000483 (S[222],C[223],S[483],C[483]);
  ha HA_00000484 (P[26][31],C[256],S[484],C[484]);
  ha HA_00000485 (S[256],C[257],S[485],C[485]);
  ha HA_00000486 (S[257],C[258],S[486],C[486]);
  fa FA_00000487 (C[224],S[258],C[259],S[487],C[487]);
  fa FA_00000488 (C[225],S[259],C[260],S[488],C[488]);
  fa FA_00000489 (C[226],S[260],C[261],S[489],C[489]);
  fa FA_00000490 (C[227],S[261],C[262],S[490],C[490]);
  fa FA_00000491 (C[228],S[262],C[263],S[491],C[491]);
  fa FA_00000492 (C[229],S[263],C[264],S[492],C[492]);
  fa FA_00000493 (C[230],S[264],C[265],S[493],C[493]);
  fa FA_00000494 (C[231],S[265],C[266],S[494],C[494]);
  fa FA_00000495 (C[232],S[266],C[267],S[495],C[495]);
  fa FA_00000496 (C[233],S[267],C[268],S[496],C[496]);
  fa FA_00000497 (C[234],S[268],C[269],S[497],C[497]);
  fa FA_00000498 (C[235],S[269],C[270],S[498],C[498]);
  fa FA_00000499 (C[236],S[270],C[271],S[499],C[499]);
  fa FA_00000500 (C[237],S[271],C[272],S[500],C[500]);
  fa FA_00000501 (C[238],S[272],C[273],S[501],C[501]);
  fa FA_00000502 (C[239],S[273],C[274],S[502],C[502]);
  fa FA_00000503 (C[240],S[274],C[275],S[503],C[503]);
  fa FA_00000504 (C[241],S[275],C[276],S[504],C[504]);
  fa FA_00000505 (C[242],S[276],C[277],S[505],C[505]);
  fa FA_00000506 (C[243],S[277],C[278],S[506],C[506]);
  fa FA_00000507 (C[244],S[278],C[279],S[507],C[507]);
  fa FA_00000508 (C[245],S[279],C[280],S[508],C[508]);
  fa FA_00000509 (C[246],S[280],C[281],S[509],C[509]);
  fa FA_00000510 (C[247],S[281],C[282],S[510],C[510]);
  fa FA_00000511 (C[248],S[282],C[283],S[511],C[511]);
  fa FA_00000512 (C[249],S[283],C[284],S[512],C[512]);
  fa FA_00000513 (C[250],S[284],C[285],S[513],C[513]);
  fa FA_00000514 (C[251],S[285],C[286],S[514],C[514]);
  fa FA_00000515 (C[252],S[286],C[287],S[515],C[515]);
  ha HA_00000516 (C[253],S[287],S[516],C[516]);
  ha HA_00000517 (C[254],P[24][0],S[517],C[517]);
  fa FA_00000518 (P[29][31],C[288],P[30][30],S[518],C[518]);
  fa FA_00000519 (S[288],C[289],P[30][29],S[519],C[519]);
  fa FA_00000520 (S[289],C[290],P[30][28],S[520],C[520]);
  fa FA_00000521 (S[290],C[291],P[30][27],S[521],C[521]);
  fa FA_00000522 (S[291],C[292],P[30][26],S[522],C[522]);
  fa FA_00000523 (S[292],C[293],P[30][25],S[523],C[523]);
  fa FA_00000524 (S[293],C[294],P[30][24],S[524],C[524]);
  fa FA_00000525 (S[294],C[295],P[30][23],S[525],C[525]);
  fa FA_00000526 (S[295],C[296],P[30][22],S[526],C[526]);
  fa FA_00000527 (S[296],C[297],P[30][21],S[527],C[527]);
  fa FA_00000528 (S[297],C[298],P[30][20],S[528],C[528]);
  fa FA_00000529 (S[298],C[299],P[30][19],S[529],C[529]);
  fa FA_00000530 (S[299],C[300],P[30][18],S[530],C[530]);
  fa FA_00000531 (S[300],C[301],P[30][17],S[531],C[531]);
  fa FA_00000532 (S[301],C[302],P[30][16],S[532],C[532]);
  fa FA_00000533 (S[302],C[303],P[30][15],S[533],C[533]);
  fa FA_00000534 (S[303],C[304],P[30][14],S[534],C[534]);
  fa FA_00000535 (S[304],C[305],P[30][13],S[535],C[535]);
  fa FA_00000536 (S[305],C[306],P[30][12],S[536],C[536]);
  fa FA_00000537 (S[306],C[307],P[30][11],S[537],C[537]);
  fa FA_00000538 (S[307],C[308],P[30][10],S[538],C[538]);
  fa FA_00000539 (S[308],C[309],P[30][9],S[539],C[539]);
  fa FA_00000540 (S[309],C[310],P[30][8],S[540],C[540]);
  fa FA_00000541 (S[310],C[311],P[30][7],S[541],C[541]);
  fa FA_00000542 (S[311],C[312],P[30][6],S[542],C[542]);
  fa FA_00000543 (S[312],C[313],P[30][5],S[543],C[543]);
  fa FA_00000544 (S[313],C[314],P[30][4],S[544],C[544]);
  fa FA_00000545 (S[314],C[315],P[30][3],S[545],C[545]);
  fa FA_00000546 (S[315],C[316],P[30][2],S[546],C[546]);
  fa FA_00000547 (S[316],C[317],P[30][1],S[547],C[547]);
  fa FA_00000548 (S[317],C[318],P[30][0],S[548],C[548]);
  ha HA_00000549 (S[318],C[319],S[549],C[549]);
  ha HA_00000550 (P[5][31],S[355],S[550],C[550]);
  ha HA_00000551 (S[32],S[356],S[551],C[551]);
  fa FA_00000552 (S[33],C[320],S[357],S[552],C[552]);
  fa FA_00000553 (S[320],C[321],S[358],S[553],C[553]);
  fa FA_00000554 (S[321],C[322],S[359],S[554],C[554]);
  fa FA_00000555 (S[322],C[323],S[360],S[555],C[555]);
  fa FA_00000556 (S[323],C[324],S[361],S[556],C[556]);
  fa FA_00000557 (S[324],C[325],S[362],S[557],C[557]);
  fa FA_00000558 (S[325],C[326],S[363],S[558],C[558]);
  fa FA_00000559 (S[326],C[327],S[364],S[559],C[559]);
  fa FA_00000560 (S[327],C[328],S[365],S[560],C[560]);
  fa FA_00000561 (S[328],C[329],S[366],S[561],C[561]);
  fa FA_00000562 (S[329],C[330],S[367],S[562],C[562]);
  fa FA_00000563 (S[330],C[331],S[368],S[563],C[563]);
  fa FA_00000564 (S[331],C[332],S[369],S[564],C[564]);
  fa FA_00000565 (S[332],C[333],S[370],S[565],C[565]);
  fa FA_00000566 (S[333],C[334],S[371],S[566],C[566]);
  fa FA_00000567 (S[334],C[335],S[372],S[567],C[567]);
  fa FA_00000568 (S[335],C[336],S[373],S[568],C[568]);
  fa FA_00000569 (S[336],C[337],S[374],S[569],C[569]);
  fa FA_00000570 (S[337],C[338],S[375],S[570],C[570]);
  fa FA_00000571 (S[338],C[339],S[376],S[571],C[571]);
  fa FA_00000572 (S[339],C[340],S[377],S[572],C[572]);
  fa FA_00000573 (S[340],C[341],S[378],S[573],C[573]);
  fa FA_00000574 (S[341],C[342],S[379],S[574],C[574]);
  fa FA_00000575 (S[342],C[343],S[380],S[575],C[575]);
  fa FA_00000576 (S[343],C[344],S[381],S[576],C[576]);
  fa FA_00000577 (S[344],C[345],S[382],S[577],C[577]);
  fa FA_00000578 (S[345],C[346],S[383],S[578],C[578]);
  fa FA_00000579 (S[346],C[347],S[384],S[579],C[579]);
  fa FA_00000580 (S[347],C[348],S[385],S[580],C[580]);
  fa FA_00000581 (S[348],C[349],C[63],S[581],C[581]);
  ha HA_00000582 (S[349],C[350],S[582],C[582]);
  ha HA_00000583 (S[350],C[351],S[583],C[583]);
  ha HA_00000584 (S[129],C[386],S[584],C[584]);
  ha HA_00000585 (S[386],C[387],S[585],C[585]);
  ha HA_00000586 (S[387],C[388],S[586],C[586]);
  fa FA_00000587 (C[352],S[388],C[389],S[587],C[587]);
  fa FA_00000588 (C[353],S[389],C[390],S[588],C[588]);
  fa FA_00000589 (C[354],S[390],C[391],S[589],C[589]);
  fa FA_00000590 (C[355],S[391],C[392],S[590],C[590]);
  fa FA_00000591 (C[356],S[392],C[393],S[591],C[591]);
  fa FA_00000592 (C[357],S[393],C[394],S[592],C[592]);
  fa FA_00000593 (C[358],S[394],C[395],S[593],C[593]);
  fa FA_00000594 (C[359],S[395],C[396],S[594],C[594]);
  fa FA_00000595 (C[360],S[396],C[397],S[595],C[595]);
  fa FA_00000596 (C[361],S[397],C[398],S[596],C[596]);
  fa FA_00000597 (C[362],S[398],C[399],S[597],C[597]);
  fa FA_00000598 (C[363],S[399],C[400],S[598],C[598]);
  fa FA_00000599 (C[364],S[400],C[401],S[599],C[599]);
  fa FA_00000600 (C[365],S[401],C[402],S[600],C[600]);
  fa FA_00000601 (C[366],S[402],C[403],S[601],C[601]);
  fa FA_00000602 (C[367],S[403],C[404],S[602],C[602]);
  fa FA_00000603 (C[368],S[404],C[405],S[603],C[603]);
  fa FA_00000604 (C[369],S[405],C[406],S[604],C[604]);
  fa FA_00000605 (C[370],S[406],C[407],S[605],C[605]);
  fa FA_00000606 (C[371],S[407],C[408],S[606],C[606]);
  fa FA_00000607 (C[372],S[408],C[409],S[607],C[607]);
  fa FA_00000608 (C[373],S[409],C[410],S[608],C[608]);
  fa FA_00000609 (C[374],S[410],C[411],S[609],C[609]);
  fa FA_00000610 (C[375],S[411],C[412],S[610],C[610]);
  fa FA_00000611 (C[376],S[412],C[413],S[611],C[611]);
  fa FA_00000612 (C[377],S[413],C[414],S[612],C[612]);
  fa FA_00000613 (C[378],S[414],C[415],S[613],C[613]);
  fa FA_00000614 (C[379],S[415],C[416],S[614],C[614]);
  fa FA_00000615 (C[380],S[416],C[417],S[615],C[615]);
  ha HA_00000616 (C[381],S[417],S[616],C[616]);
  ha HA_00000617 (C[382],S[127],S[617],C[617]);
  ha HA_00000618 (C[383],P[9][0],S[618],C[618]);
  ha HA_00000619 (C[418],S[454],S[619],C[619]);
  fa FA_00000620 (S[418],C[419],S[455],S[620],C[620]);
  fa FA_00000621 (S[419],C[420],S[456],S[621],C[621]);
  fa FA_00000622 (S[420],C[421],S[457],S[622],C[622]);
  fa FA_00000623 (S[421],C[422],S[458],S[623],C[623]);
  fa FA_00000624 (S[422],C[423],S[459],S[624],C[624]);
  fa FA_00000625 (S[423],C[424],S[460],S[625],C[625]);
  fa FA_00000626 (S[424],C[425],S[461],S[626],C[626]);
  fa FA_00000627 (S[425],C[426],S[462],S[627],C[627]);
  fa FA_00000628 (S[426],C[427],S[463],S[628],C[628]);
  fa FA_00000629 (S[427],C[428],S[464],S[629],C[629]);
  fa FA_00000630 (S[428],C[429],S[465],S[630],C[630]);
  fa FA_00000631 (S[429],C[430],S[466],S[631],C[631]);
  fa FA_00000632 (S[430],C[431],S[467],S[632],C[632]);
  fa FA_00000633 (S[431],C[432],S[468],S[633],C[633]);
  fa FA_00000634 (S[432],C[433],S[469],S[634],C[634]);
  fa FA_00000635 (S[433],C[434],S[470],S[635],C[635]);
  fa FA_00000636 (S[434],C[435],S[471],S[636],C[636]);
  fa FA_00000637 (S[435],C[436],S[472],S[637],C[637]);
  fa FA_00000638 (S[436],C[437],S[473],S[638],C[638]);
  fa FA_00000639 (S[437],C[438],S[474],S[639],C[639]);
  fa FA_00000640 (S[438],C[439],S[475],S[640],C[640]);
  fa FA_00000641 (S[439],C[440],S[476],S[641],C[641]);
  fa FA_00000642 (S[440],C[441],S[477],S[642],C[642]);
  fa FA_00000643 (S[441],C[442],S[478],S[643],C[643]);
  fa FA_00000644 (S[442],C[443],S[479],S[644],C[644]);
  fa FA_00000645 (S[443],C[444],S[480],S[645],C[645]);
  fa FA_00000646 (S[444],C[445],S[481],S[646],C[646]);
  fa FA_00000647 (S[445],C[446],S[482],S[647],C[647]);
  fa FA_00000648 (S[446],C[447],S[483],S[648],C[648]);
  fa FA_00000649 (S[447],C[448],S[223],S[649],C[649]);
  fa FA_00000650 (S[448],C[449],P[18][0],S[650],C[650]);
  ha HA_00000651 (S[449],C[450],S[651],C[651]);
  ha HA_00000652 (S[450],C[451],S[652],C[652]);
  ha HA_00000653 (S[484],C[485],S[653],C[653]);
  ha HA_00000654 (S[485],C[486],S[654],C[654]);
  ha HA_00000655 (S[486],C[487],S[655],C[655]);
  fa FA_00000656 (P[23][31],S[487],C[488],S[656],C[656]);
  fa FA_00000657 (S[224],S[488],C[489],S[657],C[657]);
  fa FA_00000658 (C[452],S[489],C[490],S[658],C[658]);
  fa FA_00000659 (C[453],S[490],C[491],S[659],C[659]);
  fa FA_00000660 (C[454],S[491],C[492],S[660],C[660]);
  fa FA_00000661 (C[455],S[492],C[493],S[661],C[661]);
  fa FA_00000662 (C[456],S[493],C[494],S[662],C[662]);
  fa FA_00000663 (C[457],S[494],C[495],S[663],C[663]);
  fa FA_00000664 (C[458],S[495],C[496],S[664],C[664]);
  fa FA_00000665 (C[459],S[496],C[497],S[665],C[665]);
  fa FA_00000666 (C[460],S[497],C[498],S[666],C[666]);
  fa FA_00000667 (C[461],S[498],C[499],S[667],C[667]);
  fa FA_00000668 (C[462],S[499],C[500],S[668],C[668]);
  fa FA_00000669 (C[463],S[500],C[501],S[669],C[669]);
  fa FA_00000670 (C[464],S[501],C[502],S[670],C[670]);
  fa FA_00000671 (C[465],S[502],C[503],S[671],C[671]);
  fa FA_00000672 (C[466],S[503],C[504],S[672],C[672]);
  fa FA_00000673 (C[467],S[504],C[505],S[673],C[673]);
  fa FA_00000674 (C[468],S[505],C[506],S[674],C[674]);
  fa FA_00000675 (C[469],S[506],C[507],S[675],C[675]);
  fa FA_00000676 (C[470],S[507],C[508],S[676],C[676]);
  fa FA_00000677 (C[471],S[508],C[509],S[677],C[677]);
  fa FA_00000678 (C[472],S[509],C[510],S[678],C[678]);
  fa FA_00000679 (C[473],S[510],C[511],S[679],C[679]);
  fa FA_00000680 (C[474],S[511],C[512],S[680],C[680]);
  fa FA_00000681 (C[475],S[512],C[513],S[681],C[681]);
  fa FA_00000682 (C[476],S[513],C[514],S[682],C[682]);
  fa FA_00000683 (C[477],S[514],C[515],S[683],C[683]);
  fa FA_00000684 (C[478],S[515],C[516],S[684],C[684]);
  fa FA_00000685 (C[479],S[516],C[517],S[685],C[685]);
  ha HA_00000686 (C[480],S[517],S[686],C[686]);
  ha HA_00000687 (C[481],C[255],S[687],C[687]);
  fa FA_00000688 (P[30][31],C[518],P[31][30],S[688],C[688]);
  fa FA_00000689 (S[518],C[519],P[31][29],S[689],C[689]);
  fa FA_00000690 (S[519],C[520],P[31][28],S[690],C[690]);
  fa FA_00000691 (S[520],C[521],P[31][27],S[691],C[691]);
  fa FA_00000692 (S[521],C[522],P[31][26],S[692],C[692]);
  fa FA_00000693 (S[522],C[523],P[31][25],S[693],C[693]);
  fa FA_00000694 (S[523],C[524],P[31][24],S[694],C[694]);
  fa FA_00000695 (S[524],C[525],P[31][23],S[695],C[695]);
  fa FA_00000696 (S[525],C[526],P[31][22],S[696],C[696]);
  fa FA_00000697 (S[526],C[527],P[31][21],S[697],C[697]);
  fa FA_00000698 (S[527],C[528],P[31][20],S[698],C[698]);
  fa FA_00000699 (S[528],C[529],P[31][19],S[699],C[699]);
  fa FA_00000700 (S[529],C[530],P[31][18],S[700],C[700]);
  fa FA_00000701 (S[530],C[531],P[31][17],S[701],C[701]);
  fa FA_00000702 (S[531],C[532],P[31][16],S[702],C[702]);
  fa FA_00000703 (S[532],C[533],P[31][15],S[703],C[703]);
  fa FA_00000704 (S[533],C[534],P[31][14],S[704],C[704]);
  fa FA_00000705 (S[534],C[535],P[31][13],S[705],C[705]);
  fa FA_00000706 (S[535],C[536],P[31][12],S[706],C[706]);
  fa FA_00000707 (S[536],C[537],P[31][11],S[707],C[707]);
  fa FA_00000708 (S[537],C[538],P[31][10],S[708],C[708]);
  fa FA_00000709 (S[538],C[539],P[31][9],S[709],C[709]);
  fa FA_00000710 (S[539],C[540],P[31][8],S[710],C[710]);
  fa FA_00000711 (S[540],C[541],P[31][7],S[711],C[711]);
  fa FA_00000712 (S[541],C[542],P[31][6],S[712],C[712]);
  fa FA_00000713 (S[542],C[543],P[31][5],S[713],C[713]);
  fa FA_00000714 (S[543],C[544],P[31][4],S[714],C[714]);
  fa FA_00000715 (S[544],C[545],P[31][3],S[715],C[715]);
  fa FA_00000716 (S[545],C[546],P[31][2],S[716],C[716]);
  fa FA_00000717 (S[546],C[547],P[31][1],S[717],C[717]);
  fa FA_00000718 (S[547],C[548],P[31][0],S[718],C[718]);
  ha HA_00000719 (S[548],C[549],S[719],C[719]);
  ha HA_00000720 (S[352],S[588],S[720],C[720]);
  ha HA_00000721 (S[353],S[589],S[721],C[721]);
  fa FA_00000722 (S[354],C[550],S[590],S[722],C[722]);
  fa FA_00000723 (S[550],C[551],S[591],S[723],C[723]);
  fa FA_00000724 (S[551],C[552],S[592],S[724],C[724]);
  fa FA_00000725 (S[552],C[553],S[593],S[725],C[725]);
  fa FA_00000726 (S[553],C[554],S[594],S[726],C[726]);
  fa FA_00000727 (S[554],C[555],S[595],S[727],C[727]);
  fa FA_00000728 (S[555],C[556],S[596],S[728],C[728]);
  fa FA_00000729 (S[556],C[557],S[597],S[729],C[729]);
  fa FA_00000730 (S[557],C[558],S[598],S[730],C[730]);
  fa FA_00000731 (S[558],C[559],S[599],S[731],C[731]);
  fa FA_00000732 (S[559],C[560],S[600],S[732],C[732]);
  fa FA_00000733 (S[560],C[561],S[601],S[733],C[733]);
  fa FA_00000734 (S[561],C[562],S[602],S[734],C[734]);
  fa FA_00000735 (S[562],C[563],S[603],S[735],C[735]);
  fa FA_00000736 (S[563],C[564],S[604],S[736],C[736]);
  fa FA_00000737 (S[564],C[565],S[605],S[737],C[737]);
  fa FA_00000738 (S[565],C[566],S[606],S[738],C[738]);
  fa FA_00000739 (S[566],C[567],S[607],S[739],C[739]);
  fa FA_00000740 (S[567],C[568],S[608],S[740],C[740]);
  fa FA_00000741 (S[568],C[569],S[609],S[741],C[741]);
  fa FA_00000742 (S[569],C[570],S[610],S[742],C[742]);
  fa FA_00000743 (S[570],C[571],S[611],S[743],C[743]);
  fa FA_00000744 (S[571],C[572],S[612],S[744],C[744]);
  fa FA_00000745 (S[572],C[573],S[613],S[745],C[745]);
  fa FA_00000746 (S[573],C[574],S[614],S[746],C[746]);
  fa FA_00000747 (S[574],C[575],S[615],S[747],C[747]);
  fa FA_00000748 (S[575],C[576],S[616],S[748],C[748]);
  fa FA_00000749 (S[576],C[577],S[617],S[749],C[749]);
  fa FA_00000750 (S[577],C[578],S[618],S[750],C[750]);
  fa FA_00000751 (S[578],C[579],C[384],S[751],C[751]);
  fa FA_00000752 (S[579],C[580],C[385],S[752],C[752]);
  ha HA_00000753 (S[580],C[581],S[753],C[753]);
  ha HA_00000754 (S[581],C[582],S[754],C[754]);
  ha HA_00000755 (S[582],C[583],S[755],C[755]);
  ha HA_00000756 (S[453],C[619],S[756],C[756]);
  ha HA_00000757 (S[619],C[620],S[757],C[757]);
  ha HA_00000758 (S[620],C[621],S[758],C[758]);
  ha HA_00000759 (S[621],C[622],S[759],C[759]);
  ha HA_00000760 (S[622],C[623],S[760],C[760]);
  fa FA_00000761 (P[14][31],S[623],C[624],S[761],C[761]);
  fa FA_00000762 (C[584],S[624],C[625],S[762],C[762]);
  fa FA_00000763 (C[585],S[625],C[626],S[763],C[763]);
  fa FA_00000764 (C[586],S[626],C[627],S[764],C[764]);
  fa FA_00000765 (C[587],S[627],C[628],S[765],C[765]);
  fa FA_00000766 (C[588],S[628],C[629],S[766],C[766]);
  fa FA_00000767 (C[589],S[629],C[630],S[767],C[767]);
  fa FA_00000768 (C[590],S[630],C[631],S[768],C[768]);
  fa FA_00000769 (C[591],S[631],C[632],S[769],C[769]);
  fa FA_00000770 (C[592],S[632],C[633],S[770],C[770]);
  fa FA_00000771 (C[593],S[633],C[634],S[771],C[771]);
  fa FA_00000772 (C[594],S[634],C[635],S[772],C[772]);
  fa FA_00000773 (C[595],S[635],C[636],S[773],C[773]);
  fa FA_00000774 (C[596],S[636],C[637],S[774],C[774]);
  fa FA_00000775 (C[597],S[637],C[638],S[775],C[775]);
  fa FA_00000776 (C[598],S[638],C[639],S[776],C[776]);
  fa FA_00000777 (C[599],S[639],C[640],S[777],C[777]);
  fa FA_00000778 (C[600],S[640],C[641],S[778],C[778]);
  fa FA_00000779 (C[601],S[641],C[642],S[779],C[779]);
  fa FA_00000780 (C[602],S[642],C[643],S[780],C[780]);
  fa FA_00000781 (C[603],S[643],C[644],S[781],C[781]);
  fa FA_00000782 (C[604],S[644],C[645],S[782],C[782]);
  fa FA_00000783 (C[605],S[645],C[646],S[783],C[783]);
  fa FA_00000784 (C[606],S[646],C[647],S[784],C[784]);
  fa FA_00000785 (C[607],S[647],C[648],S[785],C[785]);
  fa FA_00000786 (C[608],S[648],C[649],S[786],C[786]);
  fa FA_00000787 (C[609],S[649],C[650],S[787],C[787]);
  fa FA_00000788 (C[610],S[650],C[651],S[788],C[788]);
  fa FA_00000789 (C[611],S[651],C[652],S[789],C[789]);
  ha HA_00000790 (C[612],S[652],S[790],C[790]);
  ha HA_00000791 (C[613],S[451],S[791],C[791]);
  ha HA_00000792 (C[614],C[159],S[792],C[792]);
  fa FA_00000793 (C[484],C[653],S[691],S[793],C[793]);
  fa FA_00000794 (S[653],C[654],S[692],S[794],C[794]);
  fa FA_00000795 (S[654],C[655],S[693],S[795],C[795]);
  fa FA_00000796 (S[655],C[656],S[694],S[796],C[796]);
  fa FA_00000797 (S[656],C[657],S[695],S[797],C[797]);
  fa FA_00000798 (S[657],C[658],S[696],S[798],C[798]);
  fa FA_00000799 (S[658],C[659],S[697],S[799],C[799]);
  fa FA_00000800 (S[659],C[660],S[698],S[800],C[800]);
  fa FA_00000801 (S[660],C[661],S[699],S[801],C[801]);
  fa FA_00000802 (S[661],C[662],S[700],S[802],C[802]);
  fa FA_00000803 (S[662],C[663],S[701],S[803],C[803]);
  fa FA_00000804 (S[663],C[664],S[702],S[804],C[804]);
  fa FA_00000805 (S[664],C[665],S[703],S[805],C[805]);
  fa FA_00000806 (S[665],C[666],S[704],S[806],C[806]);
  fa FA_00000807 (S[666],C[667],S[705],S[807],C[807]);
  fa FA_00000808 (S[667],C[668],S[706],S[808],C[808]);
  fa FA_00000809 (S[668],C[669],S[707],S[809],C[809]);
  fa FA_00000810 (S[669],C[670],S[708],S[810],C[810]);
  fa FA_00000811 (S[670],C[671],S[709],S[811],C[811]);
  fa FA_00000812 (S[671],C[672],S[710],S[812],C[812]);
  fa FA_00000813 (S[672],C[673],S[711],S[813],C[813]);
  fa FA_00000814 (S[673],C[674],S[712],S[814],C[814]);
  fa FA_00000815 (S[674],C[675],S[713],S[815],C[815]);
  fa FA_00000816 (S[675],C[676],S[714],S[816],C[816]);
  fa FA_00000817 (S[676],C[677],S[715],S[817],C[817]);
  fa FA_00000818 (S[677],C[678],S[716],S[818],C[818]);
  fa FA_00000819 (S[678],C[679],S[717],S[819],C[819]);
  fa FA_00000820 (S[679],C[680],S[718],S[820],C[820]);
  fa FA_00000821 (S[680],C[681],S[719],S[821],C[821]);
  fa FA_00000822 (S[681],C[682],S[549],S[822],C[822]);
  fa FA_00000823 (S[682],C[683],S[319],S[823],C[823]);
  fa FA_00000824 (S[683],C[684],P[27][0],S[824],C[824]);
  ha HA_00000825 (S[684],C[685],S[825],C[825]);
  ha HA_00000826 (S[685],C[686],S[826],C[826]);
  ha HA_00000827 (S[686],C[687],S[827],C[827]);
  ha HA_00000828 (S[128],S[762],S[828],C[828]);
  ha HA_00000829 (S[584],S[763],S[829],C[829]);
  ha HA_00000830 (S[585],S[764],S[830],C[830]);
  ha HA_00000831 (S[586],S[765],S[831],C[831]);
  fa FA_00000832 (S[587],C[720],S[766],S[832],C[832]);
  fa FA_00000833 (S[720],C[721],S[767],S[833],C[833]);
  fa FA_00000834 (S[721],C[722],S[768],S[834],C[834]);
  fa FA_00000835 (S[722],C[723],S[769],S[835],C[835]);
  fa FA_00000836 (S[723],C[724],S[770],S[836],C[836]);
  fa FA_00000837 (S[724],C[725],S[771],S[837],C[837]);
  fa FA_00000838 (S[725],C[726],S[772],S[838],C[838]);
  fa FA_00000839 (S[726],C[727],S[773],S[839],C[839]);
  fa FA_00000840 (S[727],C[728],S[774],S[840],C[840]);
  fa FA_00000841 (S[728],C[729],S[775],S[841],C[841]);
  fa FA_00000842 (S[729],C[730],S[776],S[842],C[842]);
  fa FA_00000843 (S[730],C[731],S[777],S[843],C[843]);
  fa FA_00000844 (S[731],C[732],S[778],S[844],C[844]);
  fa FA_00000845 (S[732],C[733],S[779],S[845],C[845]);
  fa FA_00000846 (S[733],C[734],S[780],S[846],C[846]);
  fa FA_00000847 (S[734],C[735],S[781],S[847],C[847]);
  fa FA_00000848 (S[735],C[736],S[782],S[848],C[848]);
  fa FA_00000849 (S[736],C[737],S[783],S[849],C[849]);
  fa FA_00000850 (S[737],C[738],S[784],S[850],C[850]);
  fa FA_00000851 (S[738],C[739],S[785],S[851],C[851]);
  fa FA_00000852 (S[739],C[740],S[786],S[852],C[852]);
  fa FA_00000853 (S[740],C[741],S[787],S[853],C[853]);
  fa FA_00000854 (S[741],C[742],S[788],S[854],C[854]);
  fa FA_00000855 (S[742],C[743],S[789],S[855],C[855]);
  fa FA_00000856 (S[743],C[744],S[790],S[856],C[856]);
  fa FA_00000857 (S[744],C[745],S[791],S[857],C[857]);
  fa FA_00000858 (S[745],C[746],S[792],S[858],C[858]);
  fa FA_00000859 (S[746],C[747],C[615],S[859],C[859]);
  fa FA_00000860 (S[747],C[748],C[616],S[860],C[860]);
  fa FA_00000861 (S[748],C[749],C[617],S[861],C[861]);
  fa FA_00000862 (S[749],C[750],C[618],S[862],C[862]);
  ha HA_00000863 (S[750],C[751],S[863],C[863]);
  ha HA_00000864 (S[751],C[752],S[864],C[864]);
  ha HA_00000865 (S[752],C[753],S[865],C[865]);
  ha HA_00000866 (S[753],C[754],S[866],C[866]);
  ha HA_00000867 (S[754],C[755],S[867],C[867]);
  ha HA_00000868 (S[690],C[793],S[868],C[868]);
  ha HA_00000869 (S[793],C[794],S[869],C[869]);
  ha HA_00000870 (S[794],C[795],S[870],C[870]);
  ha HA_00000871 (S[795],C[796],S[871],C[871]);
  ha HA_00000872 (S[796],C[797],S[872],C[872]);
  ha HA_00000873 (S[797],C[798],S[873],C[873]);
  ha HA_00000874 (S[798],C[799],S[874],C[874]);
  fa FA_00000875 (S[225],S[799],C[800],S[875],C[875]);
  fa FA_00000876 (C[756],S[800],C[801],S[876],C[876]);
  fa FA_00000877 (C[757],S[801],C[802],S[877],C[877]);
  fa FA_00000878 (C[758],S[802],C[803],S[878],C[878]);
  fa FA_00000879 (C[759],S[803],C[804],S[879],C[879]);
  fa FA_00000880 (C[760],S[804],C[805],S[880],C[880]);
  fa FA_00000881 (C[761],S[805],C[806],S[881],C[881]);
  fa FA_00000882 (C[762],S[806],C[807],S[882],C[882]);
  fa FA_00000883 (C[763],S[807],C[808],S[883],C[883]);
  fa FA_00000884 (C[764],S[808],C[809],S[884],C[884]);
  fa FA_00000885 (C[765],S[809],C[810],S[885],C[885]);
  fa FA_00000886 (C[766],S[810],C[811],S[886],C[886]);
  fa FA_00000887 (C[767],S[811],C[812],S[887],C[887]);
  fa FA_00000888 (C[768],S[812],C[813],S[888],C[888]);
  fa FA_00000889 (C[769],S[813],C[814],S[889],C[889]);
  fa FA_00000890 (C[770],S[814],C[815],S[890],C[890]);
  fa FA_00000891 (C[771],S[815],C[816],S[891],C[891]);
  fa FA_00000892 (C[772],S[816],C[817],S[892],C[892]);
  fa FA_00000893 (C[773],S[817],C[818],S[893],C[893]);
  fa FA_00000894 (C[774],S[818],C[819],S[894],C[894]);
  fa FA_00000895 (C[775],S[819],C[820],S[895],C[895]);
  fa FA_00000896 (C[776],S[820],C[821],S[896],C[896]);
  fa FA_00000897 (C[777],S[821],C[822],S[897],C[897]);
  fa FA_00000898 (C[778],S[822],C[823],S[898],C[898]);
  fa FA_00000899 (C[779],S[823],C[824],S[899],C[899]);
  fa FA_00000900 (C[780],S[824],C[825],S[900],C[900]);
  fa FA_00000901 (C[781],S[825],C[826],S[901],C[901]);
  fa FA_00000902 (C[782],S[826],C[827],S[902],C[902]);
  ha HA_00000903 (C[783],S[827],S[903],C[903]);
  ha HA_00000904 (C[784],S[687],S[904],C[904]);
  ha HA_00000905 (C[785],C[482],S[905],C[905]);
  ha HA_00000906 (C[786],C[483],S[906],C[906]);
  ha HA_00000907 (S[452],S[876],S[907],C[907]);
  ha HA_00000908 (S[756],S[877],S[908],C[908]);
  ha HA_00000909 (S[757],S[878],S[909],C[909]);
  ha HA_00000910 (S[758],S[879],S[910],C[910]);
  ha HA_00000911 (S[759],S[880],S[911],C[911]);
  ha HA_00000912 (S[760],S[881],S[912],C[912]);
  fa FA_00000913 (S[761],C[828],S[882],S[913],C[913]);
  fa FA_00000914 (S[828],C[829],S[883],S[914],C[914]);
  fa FA_00000915 (S[829],C[830],S[884],S[915],C[915]);
  fa FA_00000916 (S[830],C[831],S[885],S[916],C[916]);
  fa FA_00000917 (S[831],C[832],S[886],S[917],C[917]);
  fa FA_00000918 (S[832],C[833],S[887],S[918],C[918]);
  fa FA_00000919 (S[833],C[834],S[888],S[919],C[919]);
  fa FA_00000920 (S[834],C[835],S[889],S[920],C[920]);
  fa FA_00000921 (S[835],C[836],S[890],S[921],C[921]);
  fa FA_00000922 (S[836],C[837],S[891],S[922],C[922]);
  fa FA_00000923 (S[837],C[838],S[892],S[923],C[923]);
  fa FA_00000924 (S[838],C[839],S[893],S[924],C[924]);
  fa FA_00000925 (S[839],C[840],S[894],S[925],C[925]);
  fa FA_00000926 (S[840],C[841],S[895],S[926],C[926]);
  fa FA_00000927 (S[841],C[842],S[896],S[927],C[927]);
  fa FA_00000928 (S[842],C[843],S[897],S[928],C[928]);
  fa FA_00000929 (S[843],C[844],S[898],S[929],C[929]);
  fa FA_00000930 (S[844],C[845],S[899],S[930],C[930]);
  fa FA_00000931 (S[845],C[846],S[900],S[931],C[931]);
  fa FA_00000932 (S[846],C[847],S[901],S[932],C[932]);
  fa FA_00000933 (S[847],C[848],S[902],S[933],C[933]);
  fa FA_00000934 (S[848],C[849],S[903],S[934],C[934]);
  fa FA_00000935 (S[849],C[850],S[904],S[935],C[935]);
  fa FA_00000936 (S[850],C[851],S[905],S[936],C[936]);
  fa FA_00000937 (S[851],C[852],S[906],S[937],C[937]);
  fa FA_00000938 (S[852],C[853],C[787],S[938],C[938]);
  fa FA_00000939 (S[853],C[854],C[788],S[939],C[939]);
  fa FA_00000940 (S[854],C[855],C[789],S[940],C[940]);
  fa FA_00000941 (S[855],C[856],C[790],S[941],C[941]);
  fa FA_00000942 (S[856],C[857],C[791],S[942],C[942]);
  fa FA_00000943 (S[857],C[858],C[792],S[943],C[943]);
  ha HA_00000944 (S[858],C[859],S[944],C[944]);
  ha HA_00000945 (S[859],C[860],S[945],C[945]);
  ha HA_00000946 (S[860],C[861],S[946],C[946]);
  ha HA_00000947 (S[861],C[862],S[947],C[947]);
  ha HA_00000948 (S[862],C[863],S[948],C[948]);
  ha HA_00000949 (S[863],C[864],S[949],C[949]);
  ha HA_00000950 (S[864],C[865],S[950],C[950]);
  ha HA_00000951 (S[865],C[866],S[951],C[951]);
  ha HA_00000952 (S[866],C[867],S[952],C[952]);
  ha HA_00000953 (S[689],C[868],S[953],C[953]);
  ha HA_00000954 (S[868],C[869],S[954],C[954]);
  ha HA_00000955 (S[869],C[870],S[955],C[955]);
  ha HA_00000956 (S[870],C[871],S[956],C[956]);
  ha HA_00000957 (S[871],C[872],S[957],C[957]);
  ha HA_00000958 (S[872],C[873],S[958],C[958]);
  ha HA_00000959 (S[873],C[874],S[959],C[959]);
  ha HA_00000960 (S[874],C[875],S[960],C[960]);
  fa FA_00000961 (S[875],C[907],C[876],S[961],C[961]);
  fa FA_00000962 (S[907],C[908],C[877],S[962],C[962]);
  fa FA_00000963 (S[908],C[909],C[878],S[963],C[963]);
  fa FA_00000964 (S[909],C[910],C[879],S[964],C[964]);
  fa FA_00000965 (S[910],C[911],C[880],S[965],C[965]);
  fa FA_00000966 (S[911],C[912],C[881],S[966],C[966]);
  fa FA_00000967 (S[912],C[913],C[882],S[967],C[967]);
  fa FA_00000968 (S[913],C[914],C[883],S[968],C[968]);
  fa FA_00000969 (S[914],C[915],C[884],S[969],C[969]);
  fa FA_00000970 (S[915],C[916],C[885],S[970],C[970]);
  fa FA_00000971 (S[916],C[917],C[886],S[971],C[971]);
  fa FA_00000972 (S[917],C[918],C[887],S[972],C[972]);
  fa FA_00000973 (S[918],C[919],C[888],S[973],C[973]);
  fa FA_00000974 (S[919],C[920],C[889],S[974],C[974]);
  fa FA_00000975 (S[920],C[921],C[890],S[975],C[975]);
  fa FA_00000976 (S[921],C[922],C[891],S[976],C[976]);
  fa FA_00000977 (S[922],C[923],C[892],S[977],C[977]);
  fa FA_00000978 (S[923],C[924],C[893],S[978],C[978]);
  fa FA_00000979 (S[924],C[925],C[894],S[979],C[979]);
  fa FA_00000980 (S[925],C[926],C[895],S[980],C[980]);
  fa FA_00000981 (S[926],C[927],C[896],S[981],C[981]);
  fa FA_00000982 (S[927],C[928],C[897],S[982],C[982]);
  fa FA_00000983 (S[928],C[929],C[898],S[983],C[983]);
  fa FA_00000984 (S[929],C[930],C[899],S[984],C[984]);
  fa FA_00000985 (S[930],C[931],C[900],S[985],C[985]);
  fa FA_00000986 (S[931],C[932],C[901],S[986],C[986]);
  fa FA_00000987 (S[932],C[933],C[902],S[987],C[987]);
  fa FA_00000988 (S[933],C[934],C[903],S[988],C[988]);
  fa FA_00000989 (S[934],C[935],C[904],S[989],C[989]);
  fa FA_00000990 (S[935],C[936],C[905],S[990],C[990]);
  fa FA_00000991 (S[936],C[937],C[906],S[991],C[991]);
  ha HA_00000992 (S[937],C[938],S[992],C[992]);
  ha HA_00000993 (S[938],C[939],S[993],C[993]);
  ha HA_00000994 (S[939],C[940],S[994],C[994]);
  ha HA_00000995 (S[940],C[941],S[995],C[995]);
  ha HA_00000996 (S[941],C[942],S[996],C[996]);
  ha HA_00000997 (S[942],C[943],S[997],C[997]);
  ha HA_00000998 (S[943],C[944],S[998],C[998]);
  ha HA_00000999 (S[944],C[945],S[999],C[999]);
  ha HA_00001000 (S[945],C[946],S[1000],C[1000]);
  ha HA_00001001 (S[946],C[947],S[1001],C[1001]);
  ha HA_00001002 (S[947],C[948],S[1002],C[1002]);
  ha HA_00001003 (S[948],C[949],S[1003],C[1003]);
  ha HA_00001004 (S[949],C[950],S[1004],C[1004]);
  ha HA_00001005 (S[950],C[951],S[1005],C[1005]);
  ha HA_00001006 (S[951],C[952],S[1006],C[1006]);
  ha HA_00001007 (P[31][31],C[688],S[1007],C[1007]);
  fa FA_00001008 (S[688],C[953],C[689],S[1008],C[1008]);
  fa FA_00001009 (S[953],C[954],C[690],S[1009],C[1009]);
  fa FA_00001010 (S[954],C[955],C[691],S[1010],C[1010]);
  fa FA_00001011 (S[955],C[956],C[692],S[1011],C[1011]);
  fa FA_00001012 (S[956],C[957],C[693],S[1012],C[1012]);
  fa FA_00001013 (S[957],C[958],C[694],S[1013],C[1013]);
  fa FA_00001014 (S[958],C[959],C[695],S[1014],C[1014]);
  fa FA_00001015 (S[959],C[960],C[696],S[1015],C[1015]);
  fa FA_00001016 (S[960],C[961],C[697],S[1016],C[1016]);
  fa FA_00001017 (S[961],C[962],C[698],S[1017],C[1017]);
  fa FA_00001018 (S[962],C[963],C[699],S[1018],C[1018]);
  fa FA_00001019 (S[963],C[964],C[700],S[1019],C[1019]);
  fa FA_00001020 (S[964],C[965],C[701],S[1020],C[1020]);
  fa FA_00001021 (S[965],C[966],C[702],S[1021],C[1021]);
  fa FA_00001022 (S[966],C[967],C[703],S[1022],C[1022]);
  fa FA_00001023 (S[967],C[968],C[704],S[1023],C[1023]);
  fa FA_00001024 (S[968],C[969],C[705],S[1024],C[1024]);
  fa FA_00001025 (S[969],C[970],C[706],S[1025],C[1025]);
  fa FA_00001026 (S[970],C[971],C[707],S[1026],C[1026]);
  fa FA_00001027 (S[971],C[972],C[708],S[1027],C[1027]);
  fa FA_00001028 (S[972],C[973],C[709],S[1028],C[1028]);
  fa FA_00001029 (S[973],C[974],C[710],S[1029],C[1029]);
  fa FA_00001030 (S[974],C[975],C[711],S[1030],C[1030]);
  fa FA_00001031 (S[975],C[976],C[712],S[1031],C[1031]);
  fa FA_00001032 (S[976],C[977],C[713],S[1032],C[1032]);
  fa FA_00001033 (S[977],C[978],C[714],S[1033],C[1033]);
  fa FA_00001034 (S[978],C[979],C[715],S[1034],C[1034]);
  fa FA_00001035 (S[979],C[980],C[716],S[1035],C[1035]);
  fa FA_00001036 (S[980],C[981],C[717],S[1036],C[1036]);
  fa FA_00001037 (S[981],C[982],C[718],S[1037],C[1037]);
  fa FA_00001038 (S[982],C[983],C[719],S[1038],C[1038]);
  ha HA_00001039 (S[983],C[984],S[1039],C[1039]);
  ha HA_00001040 (S[984],C[985],S[1040],C[1040]);
  ha HA_00001041 (S[985],C[986],S[1041],C[1041]);
  ha HA_00001042 (S[986],C[987],S[1042],C[1042]);
  ha HA_00001043 (S[987],C[988],S[1043],C[1043]);
  ha HA_00001044 (S[988],C[989],S[1044],C[1044]);
  ha HA_00001045 (S[989],C[990],S[1045],C[1045]);
  ha HA_00001046 (S[990],C[991],S[1046],C[1046]);
  ha HA_00001047 (S[991],C[992],S[1047],C[1047]);
  ha HA_00001048 (S[992],C[993],S[1048],C[1048]);
  ha HA_00001049 (S[993],C[994],S[1049],C[1049]);
  ha HA_00001050 (S[994],C[995],S[1050],C[1050]);
  ha HA_00001051 (S[995],C[996],S[1051],C[1051]);
  ha HA_00001052 (S[996],C[997],S[1052],C[1052]);
  ha HA_00001053 (S[997],C[998],S[1053],C[1053]);
  ha HA_00001054 (S[998],C[999],S[1054],C[1054]);
  ha HA_00001055 (S[999],C[1000],S[1055],C[1055]);
  ha HA_00001056 (S[1000],C[1001],S[1056],C[1056]);
  ha HA_00001057 (S[1001],C[1002],S[1057],C[1057]);
  ha HA_00001058 (S[1002],C[1003],S[1058],C[1058]);
  ha HA_00001059 (S[1003],C[1004],S[1059],C[1059]);
  ha HA_00001060 (S[1004],C[1005],S[1060],C[1060]);
  ha HA_00001061 (S[1005],C[1006],S[1061],C[1061]);

  assign z0[0] = P[0][0];
  assign z0[1] = S[31];
  assign z0[2] = S[351];
  assign z0[3] = S[583];
  assign z0[4] = S[755];
  assign z0[5] = S[867];
  assign z0[6] = S[952];
  assign z0[7] = S[1006];
  assign z0[8] = S[1061];
  assign z0[9] = S[1060];
  assign z0[10] = S[1059];
  assign z0[11] = S[1058];
  assign z0[12] = S[1057];
  assign z0[13] = S[1056];
  assign z0[14] = S[1055];
  assign z0[15] = S[1054];
  assign z0[16] = S[1053];
  assign z0[17] = S[1052];
  assign z0[18] = S[1051];
  assign z0[19] = S[1050];
  assign z0[20] = S[1049];
  assign z0[21] = S[1048];
  assign z0[22] = S[1047];
  assign z0[23] = S[1046];
  assign z0[24] = S[1045];
  assign z0[25] = S[1044];
  assign z0[26] = S[1043];
  assign z0[27] = S[1042];
  assign z0[28] = S[1041];
  assign z0[29] = S[1040];
  assign z0[30] = S[1039];
  assign z0[31] = S[1038];
  assign z0[32] = S[1037];
  assign z0[33] = S[1036];
  assign z0[34] = S[1035];
  assign z0[35] = S[1034];
  assign z0[36] = S[1033];
  assign z0[37] = S[1032];
  assign z0[38] = S[1031];
  assign z0[39] = S[1030];
  assign z0[40] = S[1029];
  assign z0[41] = S[1028];
  assign z0[42] = S[1027];
  assign z0[43] = S[1026];
  assign z0[44] = S[1025];
  assign z0[45] = S[1024];
  assign z0[46] = S[1023];
  assign z0[47] = S[1022];
  assign z0[48] = S[1021];
  assign z0[49] = S[1020];
  assign z0[50] = S[1019];
  assign z0[51] = S[1018];
  assign z0[52] = S[1017];
  assign z0[53] = S[1016];
  assign z0[54] = S[1015];
  assign z0[55] = S[1014];
  assign z0[56] = S[1013];
  assign z0[57] = S[1012];
  assign z0[58] = S[1011];
  assign z0[59] = S[1010];
  assign z0[60] = S[1009];
  assign z0[61] = S[1008];
  assign z0[62] = S[1007];
  assign z0[63] = 0;
  assign z1[0] = 0;
  assign z1[1] = 0;
  assign z1[2] = 0;
  assign z1[3] = 0;
  assign z1[4] = 0;
  assign z1[5] = 0;
  assign z1[6] = 0;
  assign z1[7] = 0;
  assign z1[8] = 0;
  assign z1[9] = C[1061];
  assign z1[10] = C[1060];
  assign z1[11] = C[1059];
  assign z1[12] = C[1058];
  assign z1[13] = C[1057];
  assign z1[14] = C[1056];
  assign z1[15] = C[1055];
  assign z1[16] = C[1054];
  assign z1[17] = C[1053];
  assign z1[18] = C[1052];
  assign z1[19] = C[1051];
  assign z1[20] = C[1050];
  assign z1[21] = C[1049];
  assign z1[22] = C[1048];
  assign z1[23] = C[1047];
  assign z1[24] = C[1046];
  assign z1[25] = C[1045];
  assign z1[26] = C[1044];
  assign z1[27] = C[1043];
  assign z1[28] = C[1042];
  assign z1[29] = C[1041];
  assign z1[30] = C[1040];
  assign z1[31] = C[1039];
  assign z1[32] = C[1038];
  assign z1[33] = C[1037];
  assign z1[34] = C[1036];
  assign z1[35] = C[1035];
  assign z1[36] = C[1034];
  assign z1[37] = C[1033];
  assign z1[38] = C[1032];
  assign z1[39] = C[1031];
  assign z1[40] = C[1030];
  assign z1[41] = C[1029];
  assign z1[42] = C[1028];
  assign z1[43] = C[1027];
  assign z1[44] = C[1026];
  assign z1[45] = C[1025];
  assign z1[46] = C[1024];
  assign z1[47] = C[1023];
  assign z1[48] = C[1022];
  assign z1[49] = C[1021];
  assign z1[50] = C[1020];
  assign z1[51] = C[1019];
  assign z1[52] = C[1018];
  assign z1[53] = C[1017];
  assign z1[54] = C[1016];
  assign z1[55] = C[1015];
  assign z1[56] = C[1014];
  assign z1[57] = C[1013];
  assign z1[58] = C[1012];
  assign z1[59] = C[1011];
  assign z1[60] = C[1010];
  assign z1[61] = C[1009];
  assign z1[62] = C[1008];
  assign z1[63] = C[1007];

endmodule
module ha
(
	input  [0 : 0] a,
	input  [0 : 0] b,
	output [0 : 0] s,
	output [0 : 0] c
);

	assign s = a ^ b;
	assign c = a & b;

endmodule

module fa
(
	input  [0 : 0] a,
	input  [0 : 0] b,
	input  [0 : 0] c_i,
	output [0 : 0] s,
	output [0 : 0] c_o
);

	wire s_1,c_1,c_2;

	ha ha_1_comp (.a (a), .b(b), .s(s_1), .c(c_1));
	ha ha_2_comp (.a (s_1), .b(c_i), .s(s), .c(c_2));

	assign c_o = c_1 | c_2;

endmodule
